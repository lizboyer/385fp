 

 module font_rom ( input [10:0]	addr, 
 output [7:0]	data 
); 
 
	parameter ADDR_WIDTH = 11; 
   parameter DATA_WIDTH =  8; 
	logic [ADDR_WIDTH-1:0] addr_reg; 
				 
	// ROM definition				 
	parameter [0:2**ADDR_WIDTH-1][DATA_WIDTH-1:0] ROM = 
{{7, 7, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 4, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 5, 4, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 5, 4, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 5, 5, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 5, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 5, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 5, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 5, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 5, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 7, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 4, 4, 4, 4, 4, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 0, 0, 0, 0, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 0, 0, 0, 0, 4, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 7, 7, 7, 7, 7, 7, 0, 0, 0, 0, 4, 4, 4, 0, 0, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 7, 7, 7, 7, 0, 0, 0, 0, 0, 4, 4, 0, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 0, 7, 7, 4, 0, 0, 0, 0, 0, 4, 4, 0, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 0, 4, 4, 4, 4, 0, 0, 0, 0, 0, 4, 4, 0, 4, 4, 4, 0, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 0, 4, 4, 4, 0, 0, 0, 0, 0, 0, 4, 4, 0, 0, 0, 0, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 0, 4, 4, 4, 4, 0, 0, 0, 0, 0, 4, 4, 0, 1, 1, 0, 1, 7, 7, 7, 7, 7, 7, 0, 0, 7},
{7, 7, 7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 0, 4, 4, 4, 4, 0, 0, 0, 0, 0, 4, 4, 4, 1, 1, 1, 1, 7, 7, 7, 7, 7, 0, 0, 1, 0},
{7, 7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 0, 4, 4, 4, 4, 0, 0, 0, 0, 0, 4, 4, 4, 1, 1, 0, 0, 4, 1, 1, 1, 0, 0, 0, 0, 1},
{7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 5, 5, 5, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 0, 4, 4, 4, 0, 0, 0, 0, 0, 0, 4, 4, 4, 4, 0, 4, 4, 1, 1, 1, 1, 0, 0, 0, 0, 0},
{7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 5, 5, 5, 5, 5, 5, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 0, 4, 4, 4, 0, 0, 0, 0, 0, 0, 4, 4, 4, 0, 4, 1, 1, 1, 1, 0, 1, 1, 0, 0, 0, 7},
{7, 4, 4, 4, 4, 4, 4, 4, 7, 7, 7, 5, 5, 5, 5, 5, 5, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 0, 4, 4, 4, 0, 0, 0, 0, 0, 0, 4, 4, 4, 4, 4, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 7},
{7, 4, 4, 4, 4, 4, 7, 7, 7, 7, 7, 5, 5, 5, 5, 5, 7, 5, 5, 4, 4, 5, 4, 4, 4, 4, 4, 4, 4, 5, 0, 4, 4, 0, 0, 0, 0, 0, 0, 4, 4, 4, 4, 1, 1, 1, 0, 1, 1, 0, 1, 1, 1, 1, 7},
{7, 4, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 5, 5, 5, 5, 7, 7, 5, 5, 4, 5, 4, 4, 4, 4, 4, 4, 4, 5, 0, 4, 4, 0, 0, 0, 0, 0, 0, 4, 4, 4, 4, 1, 1, 1, 1, 1, 1, 1, 1, 0, 1, 1, 7},
{7, 4, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 5, 5, 5, 7, 7, 7, 7, 5, 5, 5, 5, 4, 4, 4, 4, 4, 4, 4, 0, 4, 4, 0, 0, 0, 0, 0, 0, 4, 4, 4, 1, 1, 1, 1, 1, 0, 1, 1, 1, 1, 1, 7, 7},
{7, 4, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 5, 5, 5, 5, 7, 7, 7, 7, 7, 5, 5, 4, 4, 4, 4, 4, 4, 4, 7, 7, 7, 0, 0, 0, 0, 0, 0, 4, 4, 4, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 7, 7},
{4, 4, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 5, 5, 5, 5, 5, 7, 7, 7, 7, 5, 5, 5, 4, 4, 4, 4, 4, 4, 4, 7, 7, 7, 0, 0, 0, 0, 0, 4, 4, 4, 1, 1, 0, 0, 1, 1, 1, 1, 1, 1, 7, 7, 7},
{4, 4, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 5, 5, 5, 5, 5, 5, 5, 7, 7, 5, 5, 5, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 0, 0, 7, 4, 4, 1, 1, 0, 0, 0, 1, 1, 1, 1, 7, 7, 7, 7},
{4, 4, 0, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 5, 5, 5, 5, 0, 5, 5, 7, 5, 5, 5, 5, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 7, 7, 7, 4, 1, 1, 0, 0, 1, 1, 7, 7, 7, 7, 7, 7, 7},
{0, 0, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 5, 5, 5, 5, 5, 0, 5, 7, 5, 5, 5, 5, 5, 5, 4, 4, 4, 4, 4, 4, 4, 4, 0, 4, 4, 4, 7, 7, 7, 1, 1, 1, 1, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 0, 0, 0, 0, 5, 5, 5, 5, 0, 5, 7, 7, 7, 0, 0, 5, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 0, 4, 4, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 7, 7},
{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 4, 4, 4, 4, 0, 4, 4, 7, 0, 0, 0, 0, 0, 0, 7, 7, 7, 7, 7, 7, 7, 7, 7}
};

 
 //code 0x1 
{{7, 7, 7, 7, 7, 7, 7, 7, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 5, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 5, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 7, 5, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 7, 5, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 4, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 4, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 4, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 4, 4, 4, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 0, 0, 0, 0, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 0, 0, 0, 0, 4, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 7, 7, 7, 7, 7, 7, 0, 0, 0, 0, 4, 4, 4, 0, 0, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 7, 7, 7, 7, 0, 0, 0, 0, 0, 4, 4, 0, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 0, 7, 7, 4, 0, 0, 0, 0, 0, 4, 4, 0, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 0, 4, 4, 4, 4, 0, 0, 0, 0, 0, 4, 4, 0, 4, 4, 4, 0, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 0, 4, 4, 4, 0, 0, 0, 0, 0, 0, 4, 4, 0, 0, 0, 0, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 0, 4, 4, 4, 4, 0, 0, 0, 0, 0, 4, 4, 0, 1, 1, 0, 1, 7, 7, 7, 7, 7, 7, 0, 0, 7},
{7, 4, 4, 4, 4, 4, 4, 4, 5, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 0, 4, 4, 4, 4, 0, 0, 0, 0, 0, 4, 4, 4, 1, 1, 1, 1, 7, 7, 7, 7, 7, 0, 0, 1, 0},
{4, 4, 4, 4, 4, 4, 5, 5, 5, 5, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 0, 4, 4, 4, 4, 0, 0, 0, 0, 0, 4, 4, 4, 1, 1, 0, 0, 4, 1, 1, 1, 0, 0, 0, 0, 1},
{4, 4, 4, 4, 4, 4, 5, 5, 5, 7, 5, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 0, 4, 4, 4, 0, 0, 0, 0, 0, 0, 4, 4, 4, 4, 0, 4, 4, 1, 1, 1, 1, 0, 0, 0, 0, 0},
{4, 4, 4, 4, 4, 4, 4, 7, 7, 7, 7, 5, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 0, 4, 4, 4, 0, 0, 0, 0, 0, 0, 4, 4, 4, 0, 4, 1, 1, 1, 1, 0, 1, 1, 0, 0, 0, 7},
{7, 4, 4, 4, 4, 4, 4, 4, 7, 7, 7, 7, 5, 5, 4, 4, 4, 5, 4, 4, 4, 4, 4, 4, 4, 0, 4, 4, 4, 0, 0, 0, 0, 0, 0, 4, 4, 4, 4, 4, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 7},
{7, 7, 4, 4, 4, 4, 4, 4, 7, 7, 7, 7, 7, 5, 5, 4, 4, 5, 4, 4, 4, 4, 4, 4, 4, 4, 0, 4, 4, 0, 0, 0, 0, 0, 0, 4, 4, 4, 4, 1, 1, 1, 0, 1, 1, 0, 1, 1, 1, 1, 7},
{7, 7, 5, 5, 4, 4, 4, 4, 4, 7, 7, 7, 7, 7, 5, 5, 4, 5, 4, 4, 4, 4, 4, 4, 5, 4, 0, 4, 4, 0, 0, 0, 0, 0, 0, 4, 4, 4, 4, 1, 1, 1, 1, 1, 1, 1, 1, 0, 1, 1, 7},
{7, 7, 7, 5, 4, 4, 4, 4, 4, 7, 7, 7, 7, 7, 7, 5, 5, 5, 4, 4, 4, 4, 4, 4, 5, 4, 0, 4, 4, 0, 0, 0, 0, 0, 0, 4, 4, 4, 1, 1, 1, 1, 1, 0, 1, 1, 1, 1, 1, 7, 7},
{7, 7, 7, 5, 5, 4, 4, 0, 4, 7, 7, 7, 7, 7, 7, 7, 7, 5, 5, 4, 4, 4, 4, 4, 5, 5, 5, 5, 5, 0, 0, 0, 0, 0, 0, 4, 4, 4, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 7, 7},
{7, 7, 7, 5, 5, 4, 4, 0, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 5, 4, 4, 4, 4, 4, 4, 5, 5, 5, 5, 5, 0, 0, 0, 0, 0, 4, 4, 4, 1, 1, 0, 0, 1, 1, 1, 1, 1, 1, 7, 7, 7},
{7, 7, 7, 7, 5, 4, 0, 4, 4, 5, 5, 7, 7, 7, 7, 7, 7, 7, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 0, 0, 0, 0, 0, 7, 4, 4, 1, 1, 0, 0, 0, 1, 1, 1, 1, 7, 7, 7, 7},
{7, 7, 7, 7, 5, 5, 4, 4, 5, 0, 5, 5, 7, 7, 7, 7, 7, 7, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 0, 0, 0, 7, 7, 7, 4, 1, 1, 0, 0, 1, 1, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 5, 5, 5, 5, 5, 0, 5, 7, 7, 7, 7, 7, 7, 7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 0, 4, 4, 7, 7, 7, 7, 7, 7, 1, 1, 1, 1, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 0, 0, 5, 5, 5, 5, 5, 0, 5, 7, 7, 7, 7, 0, 0, 0, 0, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 7, 7},
{7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 4, 4, 4, 4, 4, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 7, 7, 7, 7, 7, 7, 7, 7}
};

 
 //code 0x2 
{{4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{4, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{5, 4, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 5, 4, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 5, 5, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 5, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 5, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 5, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 5, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 5, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 4, 4, 4, 4, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 0, 0, 0, 0, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 0, 0, 0, 0, 4, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 7, 7, 7, 7, 7, 7, 0, 0, 0, 0, 4, 4, 4, 0, 0, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 7, 7, 7, 7, 0, 0, 0, 0, 0, 4, 4, 0, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 0, 7, 7, 4, 0, 0, 0, 0, 0, 4, 4, 0, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 0, 4, 4, 4, 4, 0, 0, 0, 0, 0, 4, 4, 0, 4, 4, 4, 0, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 0, 4, 4, 4, 0, 0, 0, 0, 0, 0, 4, 4, 0, 0, 0, 0, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 0, 4, 4, 4, 4, 0, 0, 0, 0, 0, 4, 4, 0, 1, 1, 0, 1, 7, 7, 7, 7, 7, 7, 0, 0, 7},
{7, 7, 7, 5, 5, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 0, 4, 4, 4, 4, 0, 0, 0, 0, 0, 4, 4, 4, 1, 1, 1, 1, 7, 7, 7, 7, 7, 0, 0, 1, 0},
{7, 7, 7, 5, 5, 5, 5, 4, 4, 4, 4, 4, 4, 4, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 0, 4, 4, 4, 4, 0, 0, 0, 0, 0, 4, 4, 4, 1, 1, 0, 0, 4, 1, 1, 1, 0, 0, 0, 0, 1},
{7, 7, 7, 5, 5, 5, 5, 4, 4, 4, 4, 4, 4, 5, 4, 4, 4, 4, 4, 4, 5, 4, 4, 4, 4, 4, 4, 0, 4, 4, 4, 0, 0, 0, 0, 0, 0, 4, 4, 4, 4, 0, 4, 4, 1, 1, 1, 1, 0, 0, 0, 0, 0},
{7, 7, 7, 5, 5, 5, 5, 4, 4, 4, 4, 4, 4, 5, 4, 4, 4, 4, 4, 4, 5, 4, 4, 4, 4, 4, 4, 0, 4, 4, 4, 0, 0, 0, 0, 0, 0, 4, 4, 4, 0, 4, 1, 1, 1, 1, 0, 1, 1, 0, 0, 0, 7},
{7, 7, 7, 5, 5, 5, 5, 4, 4, 4, 4, 4, 7, 5, 5, 5, 4, 4, 4, 4, 5, 4, 4, 4, 4, 4, 4, 0, 4, 4, 4, 0, 0, 0, 0, 0, 0, 4, 4, 4, 4, 4, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 7},
{7, 7, 7, 5, 5, 5, 7, 4, 4, 4, 4, 4, 7, 7, 7, 5, 5, 4, 4, 5, 4, 4, 4, 4, 4, 5, 4, 4, 0, 4, 4, 0, 0, 0, 0, 0, 0, 4, 4, 4, 4, 1, 1, 1, 0, 1, 1, 0, 1, 1, 1, 1, 7},
{7, 7, 7, 5, 5, 5, 7, 7, 4, 4, 4, 4, 4, 7, 7, 7, 5, 5, 4, 5, 4, 4, 4, 4, 4, 5, 4, 4, 0, 4, 4, 0, 0, 0, 0, 0, 0, 4, 4, 4, 4, 1, 1, 1, 1, 1, 1, 1, 1, 0, 1, 1, 7},
{7, 7, 5, 5, 5, 5, 7, 7, 4, 4, 4, 4, 4, 7, 7, 7, 7, 5, 5, 5, 4, 4, 4, 4, 4, 5, 4, 4, 0, 4, 4, 0, 0, 0, 0, 0, 0, 4, 4, 4, 1, 1, 1, 1, 1, 0, 1, 1, 1, 1, 1, 7, 7},
{7, 5, 5, 5, 5, 5, 7, 7, 7, 4, 4, 4, 4, 7, 7, 7, 7, 7, 7, 4, 4, 4, 4, 4, 5, 4, 4, 5, 5, 7, 7, 0, 0, 0, 0, 0, 0, 4, 4, 4, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 7, 7},
{7, 5, 5, 5, 5, 5, 7, 7, 7, 4, 4, 4, 4, 4, 7, 7, 7, 7, 7, 4, 4, 4, 4, 4, 5, 5, 5, 5, 5, 5, 7, 7, 0, 0, 0, 0, 0, 4, 4, 4, 1, 1, 0, 0, 1, 1, 1, 1, 1, 1, 7, 7, 7},
{7, 5, 5, 0, 5, 5, 7, 7, 7, 7, 4, 4, 4, 4, 7, 7, 7, 7, 7, 4, 4, 4, 4, 4, 4, 4, 5, 5, 5, 5, 5, 5, 0, 0, 0, 0, 0, 7, 4, 4, 1, 1, 0, 0, 0, 1, 1, 1, 1, 7, 7, 7, 7},
{7, 5, 0, 5, 5, 7, 7, 7, 7, 7, 4, 4, 4, 4, 4, 4, 4, 7, 7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 5, 5, 5, 0, 0, 0, 5, 5, 7, 4, 1, 1, 0, 0, 1, 1, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 5, 5, 7, 7, 7, 7, 7, 7, 7, 4, 4, 4, 4, 0, 4, 4, 7, 7, 4, 4, 4, 4, 4, 4, 4, 0, 4, 4, 0, 5, 5, 5, 5, 5, 0, 5, 7, 7, 1, 1, 1, 1, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 0, 0, 0, 4, 4, 4, 4, 4, 0, 4, 0, 0, 0, 4, 4, 4, 4, 4, 4, 4, 0, 4, 0, 5, 5, 5, 5, 5, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 7, 7},
{7, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 4, 4, 4, 0, 4, 0, 0, 0, 0, 0, 0, 4, 4, 4, 4, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 7, 7, 7, 7, 7, 7, 7, 7}
};

 
 //code 0x3 
{{7, 7, 7, 7, 7, 7, 7, 7, 7, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 7, 5, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 7, 5, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 5, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 5, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 7, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 4, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 4, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 4, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 4, 4, 4, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 0, 0, 0, 0, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 0, 0, 0, 0, 4, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 7, 7, 7, 7, 7, 7, 0, 0, 0, 0, 4, 4, 4, 0, 0, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 7, 7, 7, 7, 0, 0, 0, 0, 0, 4, 4, 0, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 0, 7, 7, 4, 0, 0, 0, 0, 0, 4, 4, 0, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 0, 4, 4, 4, 4, 0, 0, 0, 0, 0, 4, 4, 0, 4, 4, 4, 0, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 0, 4, 4, 4, 0, 0, 0, 0, 0, 0, 4, 4, 0, 0, 0, 0, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 0, 4, 4, 4, 4, 0, 0, 0, 0, 0, 4, 4, 0, 1, 1, 0, 1, 7, 7, 7, 7, 7, 7, 0, 0, 7},
{7, 7, 7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 0, 4, 4, 4, 4, 0, 0, 0, 0, 0, 4, 4, 4, 1, 1, 1, 1, 7, 7, 7, 7, 7, 0, 0, 1, 0},
{7, 7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 0, 4, 4, 4, 4, 0, 0, 0, 0, 0, 4, 4, 4, 1, 1, 0, 0, 4, 1, 1, 1, 0, 0, 0, 0, 1},
{4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 5, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 0, 4, 4, 4, 0, 0, 0, 0, 0, 0, 4, 4, 4, 4, 0, 4, 4, 1, 1, 1, 1, 0, 0, 0, 0, 0},
{4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 7, 7, 5, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 0, 4, 4, 4, 0, 0, 0, 0, 0, 0, 4, 4, 4, 0, 4, 1, 1, 1, 1, 0, 1, 1, 0, 0, 0, 7},
{4, 4, 4, 4, 4, 4, 4, 4, 5, 5, 7, 7, 7, 5, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 0, 4, 4, 4, 0, 0, 0, 0, 0, 0, 4, 4, 4, 4, 4, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 7},
{4, 4, 4, 4, 4, 4, 5, 5, 5, 5, 5, 5, 7, 7, 5, 5, 4, 4, 4, 5, 4, 4, 4, 4, 4, 5, 4, 0, 4, 4, 0, 0, 0, 0, 0, 0, 4, 4, 4, 4, 1, 1, 1, 0, 1, 1, 0, 1, 1, 1, 1, 7},
{4, 4, 4, 4, 4, 7, 5, 5, 5, 5, 5, 5, 5, 7, 7, 5, 5, 4, 4, 5, 4, 4, 4, 4, 4, 5, 5, 0, 5, 4, 4, 4, 0, 0, 0, 0, 4, 4, 4, 4, 1, 1, 1, 1, 1, 1, 1, 1, 0, 1, 1, 7},
{7, 4, 4, 4, 4, 7, 7, 7, 5, 5, 5, 0, 5, 7, 7, 7, 5, 5, 5, 5, 4, 4, 4, 4, 4, 4, 7, 7, 4, 4, 4, 4, 4, 0, 0, 0, 4, 4, 4, 1, 1, 1, 1, 1, 0, 1, 1, 1, 1, 1, 7, 7},
{7, 4, 4, 4, 4, 7, 7, 7, 7, 5, 5, 0, 5, 7, 7, 7, 7, 7, 5, 5, 4, 4, 4, 4, 4, 5, 4, 4, 4, 4, 4, 0, 4, 4, 0, 0, 4, 4, 4, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 7, 7},
{7, 4, 4, 4, 4, 7, 7, 7, 7, 7, 0, 5, 5, 7, 7, 7, 7, 7, 7, 7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 0, 4, 0, 0, 4, 4, 4, 1, 1, 0, 0, 1, 1, 1, 1, 1, 1, 7, 7, 7},
{7, 4, 4, 4, 4, 4, 7, 7, 7, 7, 5, 5, 7, 7, 7, 7, 7, 7, 7, 7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 0, 0, 0, 7, 4, 4, 1, 1, 0, 0, 0, 1, 1, 1, 1, 7, 7, 7, 7},
{7, 7, 4, 4, 4, 4, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 5, 0, 0, 0, 5, 7, 7, 4, 1, 1, 0, 0, 1, 1, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 4, 4, 4, 4, 4, 0, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 4, 4, 4, 4, 4, 4, 4, 5, 5, 5, 5, 5, 5, 5, 5, 5, 7, 7, 1, 1, 1, 1, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 4, 4, 4, 4, 4, 0, 4, 0, 0, 0, 7, 7, 7, 7, 7, 7, 0, 0, 0, 4, 4, 4, 4, 5, 5, 5, 5, 5, 5, 5, 5, 5, 0, 5, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 7, 7},
{7, 0, 0, 4, 4, 4, 4, 4, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 5, 5, 5, 5, 5, 5, 5, 0, 5, 0, 0, 0, 0, 0, 0, 7, 7, 7, 7, 7, 7, 7, 7, 7}
};

 
 //code 0x4 
{{7, 7, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 4, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 5, 4, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 5, 4, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 5, 5, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 5, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 5, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 5, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 5, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 5, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 7, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 4, 4, 4, 4, 4, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 0, 0, 0, 0, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 0, 0, 0, 0, 4, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 7, 7, 7, 7, 7, 7, 0, 0, 0, 0, 4, 4, 4, 0, 0, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 7, 7, 7, 7, 0, 0, 0, 0, 0, 4, 4, 0, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 0, 7, 7, 4, 0, 0, 0, 0, 0, 4, 4, 0, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 0, 4, 4, 4, 4, 0, 0, 0, 0, 0, 4, 4, 0, 4, 4, 4, 0, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 0, 4, 4, 4, 0, 0, 0, 0, 0, 0, 4, 4, 0, 0, 0, 0, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 0, 4, 4, 4, 4, 0, 0, 0, 0, 0, 4, 4, 0, 1, 1, 0, 1, 7, 7, 7, 7, 7, 7, 0, 0, 7},
{7, 7, 7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 0, 4, 4, 4, 4, 0, 0, 0, 0, 0, 4, 4, 4, 1, 1, 1, 1, 7, 7, 7, 7, 7, 0, 0, 1, 0},
{7, 7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 0, 4, 4, 4, 4, 0, 0, 0, 0, 0, 4, 4, 4, 1, 1, 0, 0, 4, 1, 1, 1, 0, 0, 0, 0, 1},
{7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 5, 5, 5, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 0, 4, 4, 4, 0, 0, 0, 0, 0, 0, 4, 4, 4, 4, 0, 4, 4, 1, 1, 1, 1, 0, 0, 0, 0, 0},
{7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 5, 5, 5, 5, 5, 5, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 0, 4, 4, 4, 0, 0, 0, 0, 0, 0, 4, 4, 4, 0, 4, 1, 1, 1, 1, 0, 1, 1, 0, 0, 0, 7},
{7, 4, 4, 4, 4, 4, 4, 4, 7, 7, 7, 5, 5, 5, 5, 5, 5, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 0, 4, 4, 4, 0, 0, 0, 0, 0, 0, 4, 4, 4, 4, 4, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 7},
{7, 4, 4, 4, 4, 4, 7, 7, 7, 7, 7, 5, 5, 5, 5, 5, 7, 5, 5, 4, 4, 5, 4, 4, 4, 4, 4, 4, 4, 5, 0, 4, 4, 0, 0, 0, 0, 0, 0, 4, 4, 4, 4, 1, 1, 1, 0, 1, 1, 0, 1, 1, 1, 1, 7},
{7, 4, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 5, 5, 5, 5, 7, 7, 5, 5, 4, 5, 4, 4, 4, 4, 4, 4, 4, 5, 0, 4, 4, 0, 0, 0, 0, 0, 0, 4, 4, 4, 4, 1, 1, 1, 1, 1, 1, 1, 1, 0, 1, 1, 7},
{7, 4, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 5, 5, 5, 7, 7, 7, 7, 5, 5, 5, 5, 4, 4, 4, 4, 4, 4, 4, 0, 4, 4, 0, 0, 0, 0, 0, 0, 4, 4, 4, 1, 1, 1, 1, 1, 0, 1, 1, 1, 1, 1, 7, 7},
{7, 4, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 5, 5, 5, 5, 7, 7, 7, 7, 7, 5, 5, 4, 4, 4, 4, 4, 4, 4, 7, 7, 7, 0, 0, 0, 0, 0, 0, 4, 4, 4, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 7, 7},
{4, 4, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 5, 5, 5, 5, 5, 7, 7, 7, 7, 5, 5, 5, 4, 4, 4, 4, 4, 4, 4, 7, 7, 7, 0, 0, 0, 0, 0, 4, 4, 4, 1, 1, 0, 0, 1, 1, 1, 1, 1, 1, 7, 7, 7},
{4, 4, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 5, 5, 5, 5, 5, 5, 5, 7, 7, 5, 5, 5, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 0, 0, 7, 4, 4, 1, 1, 0, 0, 0, 1, 1, 1, 1, 7, 7, 7, 7},
{4, 4, 0, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 5, 5, 5, 5, 0, 5, 5, 7, 5, 5, 5, 5, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 7, 7, 7, 4, 1, 1, 0, 0, 1, 1, 7, 7, 7, 7, 7, 7, 7},
{0, 0, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 5, 5, 5, 5, 5, 0, 5, 7, 5, 5, 5, 5, 5, 5, 4, 4, 4, 4, 4, 4, 4, 4, 0, 4, 4, 4, 7, 7, 7, 1, 1, 1, 1, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 0, 0, 0, 0, 5, 5, 5, 5, 0, 5, 7, 7, 7, 0, 0, 5, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 0, 4, 4, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 7, 7},
{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 4, 4, 4, 4, 0, 4, 4, 7, 0, 0, 0, 0, 0, 0, 7, 7, 7, 7, 7, 7, 7, 7, 7}
};

 
 //code 0x5 
{{7, 7, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 4, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 5, 4, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 5, 4, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 5, 5, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 5, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 5, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 5, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 5, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 5, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 7, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 4, 4, 4, 4, 4, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 0, 0, 0, 0, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 0, 0, 0, 0, 4, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 7, 7, 7, 7, 7, 7, 0, 0, 0, 0, 4, 4, 4, 0, 0, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 7, 7, 7, 7, 0, 0, 0, 0, 0, 4, 4, 0, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 0, 7, 7, 4, 0, 0, 0, 0, 0, 4, 4, 0, 4, 4, 4, 0, 7, 7, 7, 0, 0, 7},
{7, 7, 7, 7, 7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 0, 4, 4, 4, 4, 0, 0, 0, 0, 0, 4, 4, 0, 4, 4, 0, 7, 7, 7, 0, 0, 1, 0},
{7, 7, 7, 7, 7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 0, 4, 4, 4, 0, 0, 0, 0, 0, 0, 4, 4, 0, 0, 0, 1, 7, 7, 7, 0, 0, 0, 1},
{7, 7, 7, 7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 0, 4, 4, 4, 4, 0, 0, 0, 0, 0, 4, 4, 0, 1, 1, 0, 1, 7, 7, 1, 0, 0, 0, 0},
{7, 7, 7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 0, 4, 4, 4, 4, 0, 0, 0, 0, 0, 4, 4, 4, 1, 1, 1, 0, 7, 1, 1, 0, 0, 0, 7},
{7, 7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 0, 4, 4, 4, 4, 0, 0, 0, 0, 0, 4, 4, 4, 1, 0, 0, 4, 1, 1, 1, 1, 0, 0, 1},
{7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 5, 5, 5, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 0, 4, 4, 4, 0, 0, 0, 0, 0, 0, 4, 4, 4, 0, 4, 4, 1, 1, 0, 1, 1, 1, 1, 1},
{7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 5, 5, 5, 5, 5, 5, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 0, 4, 4, 4, 0, 0, 0, 0, 0, 0, 4, 4, 4, 0, 4, 1, 1, 1, 1, 1, 1, 1, 1, 1},
{7, 4, 4, 4, 4, 4, 4, 4, 7, 7, 7, 5, 5, 5, 5, 5, 5, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 0, 4, 4, 4, 0, 0, 0, 0, 0, 0, 4, 4, 4, 4, 1, 1, 0, 1, 1, 0, 1, 1, 0, 1},
{7, 4, 4, 4, 4, 4, 7, 7, 7, 7, 7, 5, 5, 5, 5, 5, 7, 5, 5, 4, 4, 5, 4, 4, 4, 4, 4, 4, 4, 5, 0, 4, 4, 0, 0, 0, 0, 0, 0, 4, 4, 4, 4, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1},
{7, 4, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 5, 5, 5, 5, 7, 7, 5, 5, 4, 5, 4, 4, 4, 4, 4, 4, 4, 5, 0, 4, 4, 0, 0, 0, 0, 0, 0, 4, 4, 4, 4, 1, 1, 1, 1, 1, 1, 1, 1, 1, 7},
{7, 4, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 5, 5, 5, 7, 7, 7, 7, 5, 5, 5, 5, 4, 4, 4, 4, 4, 4, 4, 0, 4, 4, 0, 0, 0, 0, 0, 0, 4, 4, 4, 1, 1, 0, 0, 1, 1, 1, 1, 1, 1, 7},
{7, 4, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 5, 5, 5, 5, 7, 7, 7, 7, 7, 5, 5, 4, 4, 4, 4, 4, 4, 4, 7, 7, 7, 0, 0, 0, 0, 0, 0, 4, 4, 4, 1, 1, 0, 1, 0, 1, 1, 1, 1, 7, 7},
{4, 4, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 5, 5, 5, 5, 5, 7, 7, 7, 7, 5, 5, 5, 4, 4, 4, 4, 4, 4, 4, 7, 7, 7, 0, 0, 0, 0, 0, 4, 4, 4, 1, 1, 0, 1, 1, 1, 1, 1, 7, 7, 7},
{4, 4, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 5, 5, 5, 5, 5, 5, 5, 7, 7, 5, 5, 5, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 0, 0, 7, 4, 4, 1, 1, 1, 1, 1, 1, 7, 7, 7, 7, 7},
{4, 4, 0, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 5, 5, 5, 5, 0, 5, 5, 7, 5, 5, 5, 5, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 7, 7, 7, 4, 1, 1, 1, 1, 7, 7, 7, 7, 7, 7, 7},
{0, 0, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 5, 5, 5, 5, 5, 0, 5, 7, 5, 5, 5, 5, 5, 5, 4, 4, 4, 4, 4, 4, 4, 4, 0, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 0, 0, 0, 0, 5, 5, 5, 5, 0, 5, 7, 7, 7, 0, 0, 5, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 0, 4, 4, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 7},
{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 4, 4, 4, 4, 0, 4, 4, 7, 0, 0, 0, 0, 0, 7, 7, 7, 7, 7, 7, 7, 7}
};

 
 //code 0x6 
{{7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 0, 0, 0, 0, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 0, 0, 0, 0, 0, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 0, 4, 4, 0, 0, 7, 7, 7, 0, 0, 0, 0, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 0, 4, 4, 5, 0, 0, 7, 7, 0, 0, 0, 0, 0, 0, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 7, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 0, 4, 4, 5, 0, 7, 7, 7, 0, 0, 0, 0, 0, 0, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 5, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 0, 4, 5, 0, 0, 7, 7, 0, 0, 0, 0, 0, 0, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 5, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 0, 4, 4, 5, 0, 0, 7, 7, 0, 0, 0, 0, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 5, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 0, 4, 4, 5, 0, 7, 7, 7, 0, 0, 0, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 5, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 0, 4, 4, 5, 0, 7, 7, 7, 0, 0, 0, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 5, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 0, 4, 4, 5, 0, 7, 7, 7, 7, 0, 4, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 5, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 0, 4, 4, 5, 0, 0, 7, 7, 7, 4, 4, 4, 4, 0, 0, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 5, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 0, 4, 5, 0, 0, 7, 7, 0, 0, 4, 4, 0, 1, 1, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 5, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 0, 5, 5, 0, 0, 0, 0, 0, 4, 4, 0, 1, 1, 1, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 5, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 0, 4, 5, 5, 5, 0, 0, 4, 4, 0, 1, 1, 1, 0, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 5, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 0, 4, 5, 0, 0, 0, 4, 4, 0, 1, 1, 0, 1, 0, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 5, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 0, 0, 0, 0, 4, 4, 4, 0, 1, 1, 0, 1, 0, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 5, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 4, 4, 4, 4, 4, 0, 1, 1, 1, 0, 1, 7, 7, 7, 7, 7, 7, 0, 0, 0, 0, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 5, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 4, 4, 4, 4, 4, 0, 1, 1, 1, 1, 1, 7, 7, 7, 7, 7, 0, 0, 0, 1, 1, 0},
{7, 7, 7, 7, 7, 7, 7, 7, 7, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 4, 4, 4, 4, 4, 0, 1, 1, 1, 1, 0, 7, 7, 1, 1, 1, 0, 0, 0, 0, 1, 0},
{7, 7, 7, 7, 7, 7, 7, 4, 4, 4, 4, 4, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 4, 4, 4, 4, 4, 4, 0, 1, 1, 0, 4, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 7},
{7, 7, 7, 7, 7, 7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 4, 4, 4, 4, 4, 4, 4, 0, 1, 0, 4, 1, 1, 1, 0, 1, 1, 1, 1, 1, 1, 1, 7},
{7, 7, 7, 7, 7, 7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 0, 4, 4, 4, 4, 4, 4, 4, 4, 0, 1, 1, 1, 1, 1, 1, 1, 0, 1, 1, 1, 1, 1, 7},
{7, 7, 7, 7, 7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 4, 0, 4, 4, 4, 4, 4, 4, 4, 0, 4, 1, 1, 1, 1, 0, 1, 1, 1, 1, 1, 1, 1, 1, 7},
{7, 7, 7, 7, 7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 7, 7, 7, 7, 7, 4, 4, 4, 0, 4, 4, 4, 4, 4, 4, 4, 4, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0, 1, 1, 1, 7},
{7, 7, 7, 7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 0, 4, 4, 4, 4, 4, 4, 4, 1, 1, 1, 1, 1, 1, 1, 1, 0, 1, 1, 1, 1, 1, 1, 7},
{7, 7, 7, 7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 0, 4, 4, 4, 4, 4, 4, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 7, 7},
{7, 7, 7, 7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 0, 4, 4, 4, 4, 4, 4, 1, 1, 0, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 7, 7, 7},
{7, 7, 7, 7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 0, 0, 4, 4, 4, 4, 1, 1, 1, 0, 0, 0, 0, 0, 7, 1, 1, 1, 1, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 0, 4, 4, 4, 4, 1, 1, 1, 0, 0, 0, 0, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 0, 4, 4, 4, 4, 1, 1, 1, 0, 0, 0, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 0, 0, 4, 4, 4, 4, 1, 1, 0, 0, 0, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 0, 4, 0, 7, 7, 1, 1, 1, 0, 0, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 0, 0, 0, 7, 7, 1, 1, 1, 4, 5, 5, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 5, 4, 4, 5, 0, 7, 7, 7, 7, 1, 1, 0, 5, 0, 5, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 5, 4, 5, 7, 7, 7, 7, 7, 7, 1, 1, 0, 5, 5, 0, 5, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 5, 5, 5, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 5, 5, 7, 7, 7, 7, 7, 7, 7, 7, 1, 1, 5, 5, 5, 0, 5, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 5, 5, 5, 5, 5, 5, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 5, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 5, 5, 5, 0, 5, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 4, 4, 4, 4, 4, 4, 4, 7, 7, 7, 5, 5, 5, 5, 5, 5, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 5, 5, 5, 0, 5, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 4, 4, 4, 4, 4, 7, 7, 7, 7, 7, 5, 5, 5, 5, 5, 7, 5, 5, 4, 4, 5, 4, 4, 4, 4, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 5, 5, 5, 5, 5, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 4, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 5, 5, 5, 5, 7, 7, 5, 5, 4, 5, 4, 4, 4, 4, 4, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 5, 5, 5, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 4, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 5, 5, 5, 7, 7, 7, 7, 5, 5, 5, 5, 4, 4, 4, 4, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 4, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 5, 5, 5, 5, 7, 7, 7, 7, 7, 5, 5, 4, 4, 4, 4, 4, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{4, 4, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 5, 5, 5, 5, 5, 7, 7, 7, 7, 5, 5, 5, 4, 4, 4, 4, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{4, 4, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 5, 5, 5, 5, 5, 5, 5, 7, 7, 5, 5, 5, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{4, 4, 0, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 5, 5, 5, 5, 0, 5, 5, 7, 5, 5, 5, 5, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{0, 0, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 5, 5, 5, 5, 5, 0, 5, 7, 5, 5, 5, 5, 5, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 0, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 0, 0, 0, 0, 5, 5, 5, 5, 0, 5, 7, 7, 7, 0, 0, 5, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 7, 7, 7, 7},
{0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 4, 4, 4, 4, 4, 0, 4, 0, 0, 0, 0, 0, 7, 7, 7, 7, 7, 7, 7, 7, 7}
};

 
 //code 0x7 
{{7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 0, 0, 0, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 0, 0, 5, 0, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 0, 0, 5, 4, 0, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 0, 0, 7, 7, 7, 7, 7, 7, 7, 0, 5, 4, 4, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 0, 0, 0, 0, 7, 7, 7, 7, 7, 7, 0, 0, 5, 4, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 0, 0, 0, 0, 0, 7, 7, 7, 7, 7, 7, 0, 5, 4, 4, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 0, 0, 0, 0, 0, 7, 7, 7, 7, 7, 7, 0, 0, 5, 4, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 0, 0, 0, 7, 7, 7, 7, 7, 7, 7, 0, 5, 4, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 0, 0, 0, 7, 7, 7, 7, 7, 7, 0, 5, 4, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 0, 0, 0, 7, 4, 4, 4, 4, 7, 0, 5, 5, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 0, 0, 4, 4, 4, 4, 4, 0, 0, 5, 0, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 0, 4, 4, 4, 4, 4, 0, 0, 0, 0, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 4, 4, 4, 4, 4, 4, 0, 0, 4, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 5, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 1, 0, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 5, 5, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 1, 0, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 5, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 0, 0, 0, 0, 0, 0, 4, 4, 4, 4, 4, 1, 1, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 5, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 0, 4, 4, 4, 4, 4, 4, 0, 0, 4, 4, 4, 1, 1, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 5, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 0, 4, 4, 1, 1, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 5, 4, 4, 4, 7, 7, 7, 7, 7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 0, 4, 1, 1, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 5, 4, 4, 4, 7, 7, 7, 7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 0, 4, 1, 1, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 5, 4, 4, 4, 4, 7, 7, 4, 5, 5, 5, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 1, 1, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 7, 5, 4, 4, 4, 5, 4, 4, 4, 4, 4, 4, 5, 5, 4, 4, 4, 4, 4, 4, 4, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 7, 5, 4, 4, 4, 4, 5, 4, 4, 4, 4, 4, 4, 4, 5, 4, 4, 4, 4, 4, 4, 4, 7, 4, 4, 4, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 5, 4, 4, 4, 4},
{7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 4, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 5, 4, 4, 4, 4},
{7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 4, 4, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 5, 4, 4, 4, 4, 4, 4, 4, 5, 4},
{7, 7, 7, 7, 7, 7, 7, 7, 7, 4, 4, 4, 4, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 5, 5, 5, 4, 4, 4, 4, 4, 5, 5},
{7, 7, 7, 7, 7, 7, 7, 7, 7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 5, 5, 5, 4, 4, 4, 5, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 5, 5, 4, 4, 4, 5, 5, 7, 5, 5, 5, 5, 7, 7, 7},
{7, 7, 7, 7, 4, 4, 4, 7, 7, 4, 4, 5, 4, 4, 4, 4, 4, 4, 4, 5, 4, 4, 5, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 5, 5, 4, 4, 7, 4, 4, 5, 4, 5, 4, 5, 4, 5, 5, 4, 4, 4, 4, 5, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 5, 5, 5, 4, 4, 7, 4, 4, 5, 5, 4, 5, 5, 4, 4, 5, 4, 5, 5, 4, 4, 5, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 5, 4, 5, 4, 4, 4, 4, 4, 5, 5, 5, 5, 5, 5, 5, 5, 4, 5, 5, 5, 4, 5, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 4, 4, 5, 4, 4, 4, 4, 4, 4, 5, 5, 5, 5, 5, 5, 5, 4, 5, 4, 5, 4, 5, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 5, 4, 5, 5, 4, 4, 4, 4, 4, 4, 4, 4, 5, 5, 5, 5, 5, 4, 5, 4, 5, 4, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 5, 5, 5, 5, 4, 4, 4, 4, 4, 4, 4, 4, 7, 7, 7, 7, 7, 4, 5, 4, 5, 4, 4, 4, 5, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 5, 5, 5, 5, 4, 5, 4, 4, 4, 4, 4, 4, 7, 7, 7, 7, 7, 5, 5, 5, 5, 4, 4, 4, 5, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 5, 5, 5, 5, 4, 4, 5, 4, 4, 4, 4, 4, 5, 7, 7, 7, 7, 7, 5, 5, 5, 5, 4, 4, 5, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 5, 5, 5, 5, 4, 4, 5, 5, 4, 4, 4, 5, 7, 7, 7, 7, 7, 7, 5, 5, 5, 5, 4, 4, 5, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 5, 5, 5, 5, 4, 7, 7, 5, 5, 5, 5, 7, 7, 7, 7, 7, 7, 7, 5, 5, 5, 5, 4, 5, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{5, 5, 5, 0, 5, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 5, 5, 5, 5, 5, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{5, 5, 0, 5, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 5, 5, 5, 5, 0, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{4, 5, 0, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 4, 0, 5, 0, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 4, 5, 0, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7}
};

 
 //code 0x8 
{{7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 0, 0, 0, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 0, 0, 0, 0, 0, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 0, 0, 0, 7, 7, 7, 7, 0, 0, 0, 0, 0, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 0, 0, 0, 0, 0, 7, 7, 7, 7, 7, 0, 0, 0, 0, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 0, 0, 0, 0, 0, 0, 0, 7, 7, 7, 7, 7, 0, 0, 0, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 0, 0, 0, 7, 7, 7, 7, 7, 0, 0, 0, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 0, 0, 4, 4, 4, 4, 4, 0, 0, 0, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 4, 4, 4, 4, 7, 0, 0, 0, 0, 0, 4, 4, 4, 0, 0, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 4, 4, 4, 7, 7, 4, 4, 4, 4, 4, 4, 4, 5, 5, 4, 4, 0, 0, 4, 4, 0, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 4, 4, 4, 4, 4, 4, 4, 4, 5, 4, 4, 4, 4, 4, 4, 4, 4, 5, 5, 4, 4, 0, 4, 0, 7, 7, 7, 7},
{7, 7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 5, 4, 4, 0, 4, 7, 7, 7, 7},
{7, 7, 4, 4, 4, 4, 4, 4, 5, 5, 5, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 0, 4, 7, 7, 7},
{7, 7, 5, 5, 4, 4, 5, 5, 7, 7, 4, 4, 5, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 0, 7, 7, 7},
{7, 7, 7, 5, 5, 5, 7, 7, 7, 4, 4, 4, 4, 4, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 0, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 5, 5, 4, 4, 4, 4, 4, 4, 4, 4, 7, 7, 7},
{7, 7, 7, 7, 4, 4, 4, 7, 7, 4, 4, 5, 4, 4, 4, 4, 4, 4, 4, 5, 4, 4, 5, 4, 4, 4, 5, 4, 4, 4, 4, 7, 7},
{7, 7, 7, 7, 5, 5, 4, 4, 7, 4, 4, 5, 4, 5, 4, 5, 4, 5, 5, 4, 4, 4, 4, 5, 4, 4, 4, 5, 4, 4, 4, 7, 7},
{7, 7, 7, 5, 5, 5, 4, 4, 7, 4, 4, 5, 5, 4, 5, 5, 4, 4, 5, 4, 5, 5, 4, 4, 5, 4, 4, 5, 4, 4, 4, 7, 7},
{7, 7, 7, 5, 4, 5, 4, 4, 4, 4, 4, 5, 5, 5, 5, 5, 5, 5, 5, 4, 5, 5, 5, 4, 5, 4, 4, 5, 4, 4, 4, 4, 7},
{7, 7, 7, 4, 4, 5, 4, 4, 4, 4, 4, 4, 5, 5, 5, 5, 5, 5, 5, 4, 5, 4, 5, 4, 5, 4, 4, 5, 5, 4, 4, 4, 4},
{7, 7, 5, 4, 5, 5, 4, 4, 4, 4, 4, 4, 4, 4, 5, 5, 5, 5, 5, 4, 5, 4, 5, 4, 4, 4, 5, 7, 5, 5, 4, 4, 4},
{7, 7, 5, 5, 5, 5, 4, 4, 4, 4, 4, 4, 4, 4, 7, 7, 7, 7, 7, 4, 5, 4, 5, 4, 4, 4, 5, 7, 7, 5, 5, 4, 5},
{7, 7, 5, 5, 5, 5, 4, 5, 4, 4, 4, 4, 4, 4, 7, 7, 7, 7, 7, 5, 5, 5, 5, 4, 4, 4, 5, 7, 7, 7, 5, 5, 7},
{7, 5, 5, 5, 5, 4, 4, 5, 4, 4, 4, 4, 4, 5, 7, 7, 7, 7, 7, 5, 5, 5, 5, 4, 4, 5, 7, 7, 7, 7, 7, 7, 7},
{7, 5, 5, 5, 5, 4, 4, 5, 5, 4, 4, 4, 5, 7, 7, 7, 7, 7, 7, 5, 5, 5, 5, 4, 4, 5, 7, 7, 7, 7, 7, 7, 7},
{7, 5, 5, 5, 5, 4, 7, 7, 5, 5, 5, 5, 7, 7, 7, 7, 7, 7, 7, 5, 5, 5, 5, 4, 5, 7, 7, 7, 7, 7, 7, 7, 7},
{5, 5, 5, 0, 5, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 5, 5, 5, 5, 5, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{5, 5, 0, 5, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 5, 5, 5, 5, 0, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{4, 5, 0, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 4, 0, 5, 0, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 4, 5, 0, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7}
};

 
 //code 0x9 
{{7, 7, 7, 7, 7, 7, 0, 0, 0, 7, 7, 7, 4, 4, 7, 7, 4, 4, 7, 7, 7, 0, 0, 0, 7, 7, 7, 7, 7, 7, 7, 7, 7, 0, 0, 0, 0, 7, 7, 7, 0, 0, 7},
{7, 7, 7, 7, 0, 0, 0, 0, 0, 0, 0, 4, 4, 4, 4, 4, 4, 4, 4, 0, 0, 0, 0, 0, 0, 7, 7, 7, 0, 0, 7, 7, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0},
{7, 7, 7, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 4, 4, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7},
{7, 7, 0, 0, 0, 0, 0, 7, 7, 0, 4, 0, 1, 1, 4, 4, 1, 1, 0, 4, 0, 7, 7, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 1, 0, 1, 1, 0, 0, 7, 7, 7},
{7, 7, 0, 0, 0, 0, 0, 7, 7, 4, 0, 1, 1, 1, 4, 4, 1, 1, 1, 0, 4, 7, 7, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 7, 7},
{7, 0, 0, 0, 0, 0, 7, 7, 7, 4, 0, 1, 1, 0, 4, 4, 0, 1, 1, 0, 4, 7, 7, 7, 0, 0, 0, 0, 0, 7, 7, 7, 0, 0, 0, 0, 0, 0, 0, 7, 0, 7, 7},
{7, 0, 0, 0, 0, 0, 7, 7, 7, 4, 0, 1, 1, 0, 4, 4, 0, 1, 1, 0, 4, 7, 7, 7, 7, 7, 0, 0, 7, 7, 7, 7, 0, 0, 0, 0, 0, 0, 7, 7, 7, 7, 7},
{7, 0, 0, 0, 0, 0, 7, 7, 7, 4, 0, 1, 1, 1, 4, 4, 1, 1, 1, 0, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 0, 0, 0, 7, 7, 7, 7, 7, 7, 7},
{7, 0, 0, 0, 0, 7, 7, 7, 7, 4, 4, 0, 1, 0, 0, 0, 0, 1, 0, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 4, 4, 4, 5, 4, 7, 7, 7, 7, 7, 7},
{7, 7, 0, 0, 0, 7, 7, 7, 1, 1, 1, 4, 0, 0, 0, 0, 0, 0, 4, 1, 1, 1, 7, 7, 7, 7, 7, 7, 7, 7, 7, 4, 4, 4, 4, 5, 4, 4, 7, 7, 7, 7, 7},
{7, 7, 0, 0, 0, 7, 7, 1, 1, 1, 1, 1, 1, 0, 1, 1, 0, 1, 1, 1, 1, 1, 1, 7, 7, 7, 7, 7, 7, 7, 4, 4, 5, 4, 4, 0, 4, 4, 7, 7, 7, 7, 7},
{7, 7, 7, 0, 0, 7, 7, 1, 0, 1, 1, 0, 1, 1, 0, 0, 1, 1, 0, 1, 1, 0, 1, 7, 7, 7, 7, 7, 7, 4, 4, 4, 4, 5, 0, 4, 4, 4, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 7, 7, 7, 7, 4, 4, 4, 4, 4, 4, 5, 4, 0, 4, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 1, 1, 1, 1, 1, 0, 1, 1, 1, 1, 0, 1, 1, 1, 1, 1, 7, 7, 7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 1, 1, 0, 1, 1, 1, 0, 0, 1, 1, 1, 0, 1, 1, 7, 7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 0, 4, 4, 0, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 4, 1, 1, 1, 1, 0, 0, 0, 0, 1, 1, 1, 1, 4, 7, 4, 4, 4, 4, 4, 4, 4, 5, 7, 0, 0, 0, 0, 0, 0, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 4, 4, 4, 4, 4, 4, 5, 7, 7, 0, 0, 0, 0, 0, 0, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 4, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 4, 0, 4, 4, 4, 4, 4, 5, 7, 7, 0, 0, 0, 0, 0, 0, 1, 0, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 4, 0, 4, 0, 0, 0, 5, 0, 5, 5, 0, 0, 0, 4, 0, 4, 4, 4, 4, 4, 5, 7, 7, 7, 0, 0, 0, 0, 0, 0, 1, 1, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 4, 4, 0, 4, 4, 0, 5, 5, 5, 0, 5, 5, 0, 4, 4, 0, 4, 4, 4, 5, 5, 7, 7, 7, 7, 0, 0, 0, 0, 0, 0, 1, 1, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 4, 4, 4, 4, 0, 4, 4, 5, 5, 5, 5, 5, 5, 4, 4, 0, 4, 4, 4, 5, 5, 7, 7, 7, 7, 0, 0, 0, 0, 1, 0, 0, 1, 1, 1, 7, 0, 7},
{7, 7, 7, 7, 4, 4, 4, 4, 4, 4, 0, 4, 4, 4, 4, 4, 4, 4, 4, 0, 4, 4, 4, 5, 5, 7, 7, 7, 7, 7, 0, 0, 0, 1, 0, 0, 1, 1, 1, 1, 7, 0, 0},
{7, 7, 7, 4, 4, 4, 4, 4, 5, 4, 4, 0, 0, 0, 0, 0, 0, 0, 0, 4, 4, 4, 5, 5, 7, 7, 7, 7, 7, 7, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 7, 0, 0},
{7, 7, 4, 4, 4, 4, 4, 5, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 5, 5, 5, 7, 7, 7, 7, 7, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, 7, 0, 0},
{7, 7, 4, 4, 4, 4, 5, 5, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 5, 5, 7, 7, 7, 7, 7, 7, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0},
{7, 4, 4, 4, 4, 5, 5, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 5, 7, 7, 7, 7, 7, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 7, 7, 0, 7},
{7, 4, 4, 4, 4, 5, 7, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 5, 7, 7, 7, 7, 7, 0, 1, 1, 7, 0, 0, 1, 1, 1, 0, 0, 7, 7, 7, 7},
{4, 4, 4, 5, 5, 5, 7, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 5, 7, 7, 7, 7, 0, 1, 7, 1, 7, 7, 0, 1, 1, 1, 7, 0, 7, 7, 7, 7},
{4, 4, 4, 4, 4, 7, 7, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 5, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 0, 0, 1, 7, 7, 7, 7, 7, 7, 7},
{4, 4, 4, 4, 4, 5, 7, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 5, 7, 7, 7, 7, 7, 7, 7, 7, 7, 0, 0, 0, 7, 7, 7, 7, 7, 7, 7, 7},
{4, 4, 4, 0, 5, 5, 7, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 5, 7, 7, 7, 7, 7, 7, 7, 7, 7, 0, 7, 0, 7, 7, 7, 7, 7, 7, 7, 7},
{4, 4, 4, 4, 0, 5, 7, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 5, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{5, 4, 4, 4, 5, 7, 7, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 5, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 5, 0, 5, 5, 7, 7, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 5, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 5, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 5, 5, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 5, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 5, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 5, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 5, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 5, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7}
};

 
 //code 0xa 
{{7, 0, 0, 7, 7, 7, 0, 0, 0, 0, 7, 7, 7, 7, 7, 7, 7, 7, 7, 0, 0, 0, 7, 7, 7, 4, 4, 7, 7, 4, 4, 7, 7, 7, 0, 0, 0, 7, 7, 7, 7, 7, 7, 7, 7, 7, 0, 0, 0, 0, 7, 7, 7, 0, 0, 7},
{0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 7, 7, 0, 0, 7, 7, 7, 0, 0, 0, 0, 0, 0, 4, 4, 4, 4, 4, 4, 4, 4, 0, 0, 0, 0, 0, 0, 7, 7, 7, 0, 0, 7, 7, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0},
{7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 4, 4, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7},
{7, 7, 7, 0, 0, 1, 1, 0, 1, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 7, 7, 0, 4, 0, 1, 1, 4, 4, 1, 1, 0, 4, 0, 7, 7, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 1, 0, 1, 1, 0, 0, 7, 7, 7},
{7, 7, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 7, 7, 4, 0, 1, 1, 1, 4, 4, 1, 1, 1, 0, 4, 7, 7, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 7, 7},
{7, 7, 0, 7, 0, 0, 0, 0, 0, 0, 0, 7, 7, 7, 0, 0, 0, 0, 0, 7, 7, 7, 4, 0, 1, 1, 0, 4, 4, 0, 1, 1, 0, 4, 7, 7, 7, 0, 0, 0, 0, 0, 7, 7, 7, 0, 0, 0, 0, 0, 0, 0, 7, 0, 7, 7},
{7, 7, 7, 7, 7, 0, 0, 0, 0, 0, 0, 7, 7, 7, 7, 0, 0, 7, 7, 7, 7, 7, 4, 0, 1, 1, 0, 4, 4, 0, 1, 1, 0, 4, 7, 7, 7, 7, 7, 0, 0, 7, 7, 7, 7, 0, 0, 0, 0, 0, 0, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 0, 0, 0, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 4, 0, 1, 1, 1, 4, 4, 1, 1, 1, 0, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 0, 0, 0, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 4, 5, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 4, 4, 0, 1, 0, 0, 0, 0, 1, 0, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 4, 4, 4, 5, 4, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 4, 4, 5, 4, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 1, 1, 1, 4, 0, 0, 0, 0, 0, 0, 4, 1, 1, 1, 7, 7, 7, 7, 7, 7, 7, 7, 7, 4, 4, 4, 4, 5, 4, 4, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 4, 4, 0, 4, 4, 5, 4, 4, 7, 7, 7, 7, 7, 7, 7, 1, 1, 1, 1, 1, 1, 0, 1, 1, 0, 1, 1, 1, 1, 1, 1, 7, 7, 7, 7, 7, 7, 7, 4, 4, 5, 4, 4, 0, 4, 4, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 4, 4, 4, 0, 5, 4, 4, 4, 4, 7, 7, 7, 7, 7, 7, 1, 0, 1, 1, 0, 1, 1, 0, 0, 1, 1, 0, 1, 1, 0, 1, 7, 7, 7, 7, 7, 7, 4, 4, 4, 4, 5, 0, 4, 4, 4, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 4, 0, 4, 5, 4, 4, 4, 4, 4, 4, 7, 7, 7, 7, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 7, 7, 7, 7, 4, 4, 4, 4, 4, 4, 5, 4, 0, 4, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 7, 7, 7, 1, 1, 1, 1, 1, 0, 1, 1, 1, 1, 0, 1, 1, 1, 1, 1, 7, 7, 7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 0, 4, 4, 0, 4, 4, 4, 4, 4, 4, 4, 4, 4, 7, 7, 1, 1, 0, 1, 1, 1, 0, 0, 1, 1, 1, 0, 1, 1, 7, 7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 0, 4, 4, 0, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 0, 0, 0, 0, 0, 0, 7, 5, 4, 4, 4, 4, 4, 4, 4, 7, 4, 1, 1, 1, 1, 0, 0, 0, 0, 1, 1, 1, 1, 4, 7, 4, 4, 4, 4, 4, 4, 4, 5, 7, 0, 0, 0, 0, 0, 0, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 0, 0, 0, 0, 0, 0, 7, 7, 5, 4, 4, 4, 4, 4, 4, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 4, 4, 4, 4, 4, 4, 5, 7, 7, 0, 0, 0, 0, 0, 0, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 0, 1, 0, 0, 0, 0, 0, 0, 7, 7, 5, 4, 4, 4, 4, 4, 0, 4, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 4, 0, 4, 4, 4, 4, 4, 5, 7, 7, 0, 0, 0, 0, 0, 0, 1, 0, 7, 7, 7, 7},
{7, 7, 7, 7, 1, 1, 0, 0, 0, 0, 0, 0, 7, 7, 7, 5, 4, 4, 4, 4, 4, 0, 4, 0, 0, 0, 5, 5, 5, 5, 0, 0, 0, 4, 0, 4, 4, 4, 4, 4, 5, 7, 7, 7, 0, 0, 0, 0, 0, 0, 1, 1, 7, 7, 7, 7},
{7, 7, 7, 7, 1, 1, 0, 0, 0, 0, 0, 0, 7, 7, 7, 7, 5, 5, 4, 4, 4, 0, 4, 4, 0, 5, 5, 0, 0, 5, 5, 0, 4, 4, 0, 4, 4, 4, 5, 5, 7, 7, 7, 7, 0, 0, 0, 0, 0, 0, 1, 1, 7, 7, 7, 7},
{7, 0, 7, 1, 1, 1, 0, 0, 1, 0, 0, 0, 0, 7, 7, 7, 7, 5, 5, 4, 4, 4, 0, 4, 4, 5, 5, 5, 5, 5, 5, 4, 4, 0, 4, 4, 4, 5, 5, 7, 7, 7, 7, 0, 0, 0, 0, 1, 0, 0, 1, 1, 1, 7, 0, 7},
{0, 0, 7, 1, 1, 1, 1, 0, 0, 1, 0, 0, 0, 7, 7, 7, 7, 7, 5, 5, 4, 4, 4, 0, 4, 4, 4, 4, 4, 4, 4, 4, 0, 4, 4, 4, 5, 5, 7, 7, 7, 7, 7, 0, 0, 0, 1, 0, 0, 1, 1, 1, 1, 7, 0, 0},
{0, 0, 7, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 7, 7, 7, 7, 7, 7, 5, 5, 4, 4, 4, 0, 0, 0, 0, 0, 0, 0, 0, 4, 4, 4, 5, 5, 7, 7, 7, 7, 7, 7, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 7, 0, 0},
{0, 0, 7, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 7, 7, 7, 7, 7, 5, 5, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 5, 5, 5, 7, 7, 7, 7, 7, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, 7, 0, 0},
{0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 7, 7, 7, 7, 7, 7, 5, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 5, 5, 7, 7, 7, 7, 7, 7, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0},
{7, 0, 7, 7, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 7, 7, 7, 7, 7, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 5, 7, 7, 7, 7, 7, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 7, 7, 0, 7},
{7, 7, 7, 7, 0, 0, 1, 1, 1, 0, 0, 7, 1, 1, 0, 7, 7, 7, 7, 7, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 5, 7, 7, 7, 7, 7, 0, 1, 1, 7, 0, 0, 1, 1, 1, 0, 0, 7, 7, 7, 7},
{7, 7, 7, 7, 0, 7, 1, 1, 1, 0, 7, 7, 1, 7, 1, 0, 7, 7, 7, 7, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 5, 7, 7, 7, 7, 0, 1, 7, 1, 7, 7, 0, 1, 1, 1, 7, 0, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 1, 0, 0, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 5, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 0, 0, 1, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 0, 0, 0, 7, 7, 7, 7, 7, 7, 7, 7, 7, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 5, 7, 7, 7, 7, 7, 7, 7, 7, 7, 0, 0, 0, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 0, 7, 0, 7, 7, 7, 7, 7, 7, 7, 7, 7, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 5, 7, 7, 7, 7, 7, 7, 7, 7, 7, 0, 7, 0, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 5, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 5, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 5, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 5, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 5, 5, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 5, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 5, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 5, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 5, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 5, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7}
};

 
 //code 0xb 
{{7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 1, 0, 0, 0, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 0, 1, 0, 0, 0, 0, 0, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 0, 0, 0, 1, 1, 0, 0, 0, 0, 0, 0, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 0, 1, 1, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 0, 0, 1, 1, 1, 0, 0, 0, 0, 1, 1, 0, 0, 0, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 0, 0, 0, 1, 1, 1, 1, 1, 0, 0, 1, 0, 0, 0, 0, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 0, 0, 1, 1, 1, 1, 1, 1, 0, 0, 1, 1, 0, 0, 0, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 0, 0, 0, 1, 1, 1, 1, 1, 1, 0, 0, 0, 1, 0, 0, 0, 0, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 0, 0, 1, 1, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 0, 0, 0, 1, 1, 1, 1, 1, 1, 1, 1, 0, 0, 0, 7, 7, 7, 0, 0, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 0, 0, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0, 0, 0, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 0, 0, 0, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 0, 0, 0, 0, 0, 1, 1, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 0, 0, 0, 1, 1, 1, 1, 1, 1, 1, 1, 0, 0, 0, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 0, 0, 7, 1, 1, 1, 1, 1, 1, 7, 0, 0, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 0, 0, 7, 7, 7, 7, 7, 7, 7, 7, 0, 0, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 0, 0, 7, 7, 7, 0, 0, 0, 0, 7, 7, 7, 7, 7, 7, 7, 7, 7, 0, 0, 0, 7, 7, 7, 4, 4, 7, 7, 4, 4, 7, 7, 7, 0, 0, 0, 7, 7, 7, 7, 7, 7, 7, 7, 7, 0, 0, 0, 0, 7, 7, 7, 0, 0, 7},
{0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 7, 7, 0, 0, 7, 7, 7, 0, 0, 0, 0, 0, 0, 4, 4, 4, 4, 4, 4, 4, 4, 0, 0, 0, 0, 0, 0, 7, 7, 7, 0, 0, 7, 7, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0},
{7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 4, 4, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7},
{7, 7, 7, 0, 0, 1, 1, 0, 1, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 7, 7, 0, 4, 0, 1, 1, 4, 4, 1, 1, 0, 4, 0, 7, 7, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 1, 0, 1, 1, 0, 0, 7, 7, 7},
{7, 7, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0, 7, 7, 4, 0, 1, 1, 1, 4, 4, 1, 1, 1, 0, 4, 7, 7, 0, 0, 0, 0, 0, 0, 0, 7, 0, 0, 0, 0, 1, 1, 0, 0, 0, 0, 7, 7},
{7, 7, 0, 7, 0, 0, 0, 0, 0, 0, 0, 7, 7, 7, 0, 0, 0, 0, 0, 7, 7, 7, 4, 0, 1, 1, 0, 4, 4, 0, 1, 1, 0, 4, 7, 7, 7, 0, 0, 0, 0, 0, 7, 7, 7, 0, 0, 0, 0, 0, 0, 0, 7, 0, 7, 7},
{7, 7, 7, 7, 7, 0, 0, 0, 0, 0, 0, 7, 7, 7, 7, 0, 0, 7, 7, 7, 7, 7, 4, 0, 1, 1, 0, 4, 4, 0, 1, 1, 0, 4, 7, 7, 7, 7, 7, 0, 0, 7, 7, 7, 7, 0, 0, 0, 0, 0, 0, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 0, 0, 0, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 4, 0, 1, 1, 1, 4, 4, 1, 1, 1, 0, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 0, 0, 0, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 4, 5, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 4, 4, 0, 1, 0, 0, 0, 0, 1, 0, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 4, 4, 4, 5, 4, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 4, 4, 5, 4, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 1, 1, 1, 4, 0, 0, 0, 0, 0, 0, 4, 1, 1, 1, 7, 7, 7, 7, 7, 7, 7, 7, 7, 4, 4, 4, 4, 5, 4, 4, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 4, 4, 0, 4, 4, 5, 4, 4, 7, 7, 7, 7, 7, 7, 7, 1, 1, 1, 1, 1, 1, 0, 1, 1, 0, 1, 1, 1, 1, 1, 1, 7, 7, 7, 7, 7, 7, 7, 4, 4, 5, 4, 4, 0, 4, 4, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 4, 4, 4, 0, 5, 4, 4, 4, 4, 7, 7, 7, 7, 7, 7, 1, 0, 1, 1, 0, 1, 1, 0, 0, 1, 1, 0, 1, 1, 0, 1, 7, 7, 7, 7, 7, 7, 4, 4, 4, 4, 5, 0, 4, 4, 4, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 4, 0, 4, 5, 4, 4, 4, 4, 4, 4, 7, 7, 7, 7, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 7, 7, 7, 7, 4, 4, 4, 4, 4, 4, 5, 4, 0, 4, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 7, 7, 7, 1, 1, 1, 1, 1, 0, 1, 1, 1, 1, 0, 1, 1, 1, 1, 1, 7, 7, 7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 0, 4, 4, 0, 4, 4, 4, 4, 4, 4, 4, 4, 4, 7, 7, 1, 1, 0, 1, 1, 1, 0, 0, 1, 1, 1, 0, 1, 1, 7, 7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 0, 4, 4, 0, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 0, 0, 0, 0, 0, 0, 7, 5, 4, 4, 4, 4, 4, 4, 4, 7, 4, 1, 1, 1, 1, 0, 0, 0, 0, 1, 1, 1, 1, 4, 7, 4, 4, 4, 4, 4, 4, 4, 5, 7, 0, 0, 0, 0, 0, 0, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 0, 0, 0, 0, 0, 0, 7, 7, 5, 4, 4, 4, 4, 4, 4, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 4, 4, 4, 4, 4, 4, 5, 7, 7, 0, 0, 0, 0, 0, 0, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 0, 1, 0, 0, 0, 0, 0, 0, 7, 7, 5, 4, 4, 4, 4, 4, 0, 4, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 4, 0, 4, 4, 4, 4, 4, 5, 7, 7, 0, 0, 0, 0, 0, 0, 1, 0, 7, 7, 7, 7},
{7, 7, 7, 7, 1, 1, 0, 0, 0, 0, 0, 0, 7, 7, 7, 5, 4, 4, 4, 4, 4, 0, 4, 0, 0, 0, 5, 5, 5, 5, 0, 0, 0, 4, 0, 4, 4, 4, 4, 4, 5, 7, 7, 7, 0, 0, 0, 0, 0, 0, 1, 1, 7, 7, 7, 7},
{7, 7, 7, 7, 1, 1, 0, 0, 0, 0, 0, 0, 7, 7, 7, 7, 5, 5, 4, 4, 4, 0, 4, 4, 0, 5, 5, 0, 0, 5, 5, 0, 4, 4, 0, 4, 4, 4, 5, 5, 7, 7, 7, 7, 0, 0, 0, 0, 0, 0, 1, 1, 7, 7, 7, 7},
{7, 0, 7, 1, 1, 1, 0, 0, 1, 0, 0, 0, 0, 7, 7, 7, 7, 5, 5, 4, 4, 4, 0, 4, 4, 5, 5, 5, 5, 5, 5, 4, 4, 0, 4, 4, 4, 5, 5, 7, 7, 7, 7, 0, 0, 0, 0, 1, 0, 0, 1, 1, 1, 7, 0, 7},
{0, 0, 7, 1, 1, 1, 1, 0, 0, 1, 0, 0, 0, 7, 7, 7, 7, 7, 5, 5, 4, 4, 4, 0, 4, 4, 4, 4, 4, 4, 4, 4, 0, 4, 4, 4, 5, 5, 7, 7, 7, 7, 7, 0, 0, 0, 1, 0, 0, 1, 1, 1, 1, 7, 0, 0},
{0, 0, 7, 1, 0, 0, 1, 0, 0, 1, 0, 0, 0, 7, 7, 7, 7, 7, 7, 5, 5, 4, 4, 4, 0, 0, 0, 0, 0, 0, 0, 0, 4, 4, 4, 5, 5, 7, 7, 7, 7, 7, 7, 0, 0, 0, 1, 0, 0, 1, 0, 0, 1, 7, 0, 0},
{0, 0, 7, 1, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 7, 7, 7, 7, 7, 5, 5, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 5, 5, 5, 7, 7, 7, 7, 7, 0, 0, 0, 1, 0, 0, 1, 0, 0, 0, 1, 7, 0, 0},
{0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 1, 1, 0, 0, 7, 7, 7, 7, 7, 7, 5, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 5, 5, 7, 7, 7, 7, 7, 7, 0, 0, 1, 1, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0},
{7, 0, 7, 7, 0, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 7, 7, 7, 7, 7, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 5, 7, 7, 7, 7, 7, 0, 0, 1, 1, 0, 0, 0, 1, 0, 0, 0, 7, 7, 0, 7},
{7, 7, 7, 7, 0, 0, 1, 1, 1, 0, 0, 7, 1, 1, 0, 7, 7, 7, 7, 7, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 5, 7, 7, 7, 7, 7, 0, 1, 1, 7, 0, 0, 1, 1, 1, 0, 0, 7, 7, 7, 7},
{7, 7, 7, 7, 0, 7, 1, 1, 1, 0, 7, 7, 1, 7, 1, 0, 7, 7, 7, 7, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 5, 7, 7, 7, 7, 0, 1, 7, 1, 7, 7, 0, 1, 1, 1, 7, 0, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 1, 0, 0, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 5, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 0, 0, 1, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 0, 0, 0, 7, 7, 7, 7, 7, 7, 7, 7, 7, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 5, 7, 7, 7, 7, 7, 7, 7, 7, 7, 0, 0, 0, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 0, 7, 0, 7, 7, 7, 7, 7, 7, 7, 7, 7, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 5, 7, 7, 7, 7, 7, 7, 7, 7, 7, 0, 7, 0, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 5, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 5, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 5, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 5, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 5, 5, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 5, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 5, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 5, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 5, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 5, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7}
};

 
 //code 0xc 
{{7, 7, 7, 7, 7, 0, 0, 0, 7, 7, 7, 4, 4, 7, 7, 4, 4, 7, 7, 7, 0, 0, 0, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 0, 0, 0, 0, 0, 0, 0, 4, 4, 4, 4, 4, 4, 4, 4, 0, 0, 0, 0, 0, 0, 7, 7, 7, 0, 0},
{7, 7, 0, 0, 0, 0, 0, 0, 0, 0, 4, 0, 0, 4, 4, 0, 0, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},
{7, 0, 0, 0, 0, 0, 7, 7, 0, 4, 0, 1, 1, 4, 4, 1, 1, 0, 4, 0, 7, 7, 0, 0, 0, 0, 0, 0, 0},
{7, 0, 0, 0, 0, 0, 7, 7, 4, 0, 1, 1, 1, 4, 4, 1, 1, 1, 0, 4, 7, 7, 0, 0, 0, 0, 0, 0, 0},
{0, 0, 0, 0, 0, 7, 7, 7, 4, 0, 1, 0, 1, 4, 4, 1, 0, 1, 0, 4, 7, 7, 7, 0, 0, 0, 0, 0, 7},
{0, 0, 0, 0, 0, 7, 7, 7, 4, 0, 1, 1, 0, 4, 4, 0, 1, 1, 0, 4, 7, 7, 7, 7, 7, 0, 0, 7, 7},
{0, 0, 0, 0, 0, 7, 7, 7, 4, 0, 1, 1, 1, 4, 4, 1, 1, 1, 0, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{0, 0, 0, 0, 7, 7, 7, 7, 4, 4, 0, 1, 0, 0, 0, 0, 1, 0, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 0, 0, 0, 7, 7, 7, 1, 1, 1, 4, 0, 0, 0, 0, 0, 0, 4, 1, 1, 1, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 0, 0, 0, 7, 7, 1, 1, 1, 1, 1, 1, 0, 1, 1, 0, 1, 1, 1, 1, 1, 1, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 0, 0, 7, 7, 1, 0, 1, 1, 0, 1, 1, 0, 0, 1, 1, 0, 1, 1, 0, 1, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 1, 1, 1, 1, 1, 0, 1, 1, 1, 1, 0, 1, 1, 1, 1, 1, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 4, 4, 0, 1, 1, 0, 1, 1, 1, 0, 0, 1, 1, 1, 0, 1, 1, 0, 4, 4, 7, 7, 7, 7, 7},
{7, 7, 7, 4, 4, 4, 1, 0, 1, 1, 1, 1, 0, 1, 1, 0, 1, 1, 1, 1, 0, 1, 4, 4, 4, 7, 7, 7, 7},
{7, 7, 4, 4, 4, 4, 1, 1, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 0, 0, 1, 1, 4, 4, 4, 4, 7, 7, 7},
{7, 7, 4, 4, 4, 4, 1, 0, 1, 1, 1, 0, 1, 1, 1, 1, 0, 1, 1, 1, 0, 1, 4, 4, 4, 4, 7, 7, 7},
{7, 4, 4, 4, 4, 0, 4, 0, 0, 1, 0, 0, 0, 1, 1, 0, 0, 0, 4, 4, 0, 0, 0, 4, 4, 4, 4, 7, 7},
{7, 4, 4, 4, 4, 0, 4, 4, 1, 1, 1, 0, 1, 1, 1, 1, 4, 4, 0, 4, 4, 0, 0, 4, 4, 4, 4, 7, 7},
{7, 4, 4, 4, 4, 0, 0, 4, 4, 1, 1, 1, 1, 1, 1, 1, 4, 4, 4, 4, 4, 0, 4, 4, 4, 4, 4, 7, 7},
{7, 5, 4, 4, 4, 4, 0, 0, 4, 4, 4, 1, 1, 1, 1, 4, 0, 4, 4, 4, 4, 0, 4, 4, 4, 4, 4, 4, 7},
{7, 5, 4, 4, 4, 4, 4, 0, 0, 0, 4, 4, 4, 4, 4, 4, 4, 0, 4, 4, 4, 4, 0, 0, 4, 4, 4, 4, 7},
{7, 5, 4, 4, 4, 4, 4, 4, 4, 0, 0, 0, 0, 0, 0, 4, 4, 4, 4, 4, 4, 4, 4, 4, 0, 4, 4, 4, 7},
{7, 7, 5, 4, 4, 4, 4, 4, 4, 4, 5, 5, 5, 4, 4, 5, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 5, 7},
{7, 7, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 5, 4, 4, 4, 5, 5, 4, 4, 4, 4, 4, 4, 4, 4, 5, 7},
{7, 7, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 5, 4, 4, 4, 4, 5, 4, 4, 4, 4, 4, 4, 5, 5, 7},
{7, 7, 7, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 0, 5, 4, 4, 4, 4, 4, 5, 4, 4, 4, 4, 4, 5, 7, 7},
{7, 7, 7, 7, 5, 5, 4, 4, 4, 4, 4, 4, 4, 4, 0, 4, 4, 4, 4, 4, 5, 5, 5, 4, 4, 5, 5, 7, 7},
{7, 7, 7, 7, 7, 7, 5, 5, 5, 4, 0, 4, 4, 4, 5, 4, 4, 4, 4, 4, 4, 5, 7, 5, 5, 5, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 5, 4, 5, 5, 4, 0, 4, 5, 4, 4, 4, 4, 4, 4, 4, 5, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 5, 4, 4, 5, 5, 5, 0, 4, 4, 4, 4, 4, 4, 4, 4, 5, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 5, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 5, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 5, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 5, 5, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 5, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 5, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 5, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 5, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 5, 7, 7, 7, 7, 7, 7, 7, 7}
};

 
 //code 0xd 
{{7, 7, 7, 7, 7, 0, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 0, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 0, 0, 0, 0, 0, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 0, 0, 0, 0, 7, 7, 7, 0, 0},
{7, 7, 0, 0, 0, 0, 0, 0, 0, 7, 7, 4, 4, 7, 7, 4, 4, 7, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},
{7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 4, 4, 4, 4, 4, 4, 4, 4, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0},
{7, 0, 0, 0, 0, 0, 7, 0, 0, 0, 4, 0, 0, 4, 4, 0, 0, 4, 0, 0, 0, 7, 0, 0, 0, 0, 0, 0, 0},
{0, 0, 0, 0, 0, 7, 7, 7, 0, 4, 0, 1, 1, 4, 4, 1, 1, 0, 4, 0, 7, 7, 7, 0, 0, 0, 0, 0, 7},
{0, 0, 0, 0, 0, 7, 7, 7, 4, 0, 1, 1, 1, 4, 4, 1, 1, 1, 0, 4, 7, 7, 7, 7, 7, 0, 0, 7, 7},
{0, 0, 0, 0, 0, 7, 7, 7, 4, 0, 1, 0, 1, 4, 4, 1, 0, 1, 0, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{0, 0, 0, 0, 7, 7, 7, 7, 4, 0, 1, 1, 0, 4, 4, 0, 1, 1, 0, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 0, 0, 0, 7, 7, 7, 7, 4, 0, 1, 1, 1, 4, 4, 1, 1, 1, 0, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 0, 0, 0, 7, 7, 7, 7, 4, 4, 0, 1, 0, 0, 0, 0, 1, 0, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 0, 0, 7, 7, 7, 1, 1, 1, 4, 0, 0, 0, 0, 0, 0, 4, 1, 1, 1, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 1, 1, 1, 1, 1, 1, 0, 1, 1, 0, 1, 1, 1, 1, 1, 1, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 1, 0, 1, 1, 0, 1, 1, 0, 0, 1, 1, 0, 1, 1, 0, 1, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 4, 4, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 4, 4, 7, 7, 7, 7, 7},
{7, 7, 7, 4, 4, 4, 1, 1, 1, 1, 1, 0, 1, 1, 1, 1, 0, 1, 1, 1, 1, 1, 4, 4, 4, 7, 7, 7, 7},
{7, 7, 4, 4, 4, 4, 0, 1, 1, 0, 1, 1, 1, 0, 0, 1, 1, 1, 0, 1, 1, 0, 4, 4, 4, 4, 7, 7, 7},
{7, 7, 4, 4, 4, 4, 1, 0, 1, 1, 1, 1, 0, 1, 1, 0, 1, 1, 1, 1, 0, 1, 4, 4, 4, 4, 7, 7, 7},
{7, 4, 4, 4, 4, 0, 1, 1, 0, 0, 0, 0, 1, 1, 1, 1, 0, 0, 4, 4, 0, 1, 0, 4, 4, 4, 4, 7, 7},
{7, 4, 4, 4, 4, 0, 4, 0, 1, 1, 1, 0, 1, 1, 1, 0, 4, 4, 0, 4, 4, 0, 0, 4, 4, 4, 4, 7, 7},
{7, 4, 4, 4, 4, 0, 4, 4, 1, 1, 1, 0, 1, 1, 1, 0, 4, 4, 4, 4, 4, 0, 4, 4, 4, 4, 4, 7, 7},
{7, 5, 4, 4, 4, 4, 0, 4, 4, 4, 1, 1, 1, 1, 1, 4, 0, 4, 4, 4, 4, 0, 4, 4, 4, 4, 4, 4, 7},
{7, 5, 4, 4, 4, 4, 4, 0, 0, 4, 4, 4, 4, 4, 4, 4, 4, 0, 4, 4, 4, 4, 0, 0, 4, 4, 4, 4, 7},
{7, 5, 4, 4, 4, 4, 4, 4, 4, 0, 0, 0, 0, 0, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 0, 4, 4, 4, 7},
{7, 7, 5, 4, 4, 4, 4, 4, 4, 4, 5, 5, 5, 4, 4, 5, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 5, 7},
{7, 7, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 5, 4, 4, 4, 5, 5, 4, 4, 4, 4, 4, 4, 4, 4, 5, 7},
{7, 7, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 5, 4, 4, 4, 4, 5, 4, 4, 4, 4, 4, 4, 5, 5, 7},
{7, 7, 7, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 0, 5, 4, 4, 4, 4, 4, 5, 4, 4, 4, 4, 4, 5, 7, 7},
{7, 7, 7, 7, 5, 5, 4, 4, 4, 4, 4, 4, 4, 4, 0, 4, 4, 4, 4, 4, 5, 5, 5, 4, 4, 5, 5, 7, 7},
{7, 7, 7, 7, 7, 7, 5, 5, 5, 4, 0, 4, 4, 4, 5, 4, 4, 4, 4, 4, 4, 5, 7, 5, 5, 5, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 5, 4, 5, 5, 4, 0, 4, 5, 4, 4, 4, 4, 4, 4, 4, 5, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 5, 4, 4, 5, 5, 5, 0, 4, 4, 4, 4, 4, 4, 4, 4, 5, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 5, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 5, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 5, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 5, 5, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 5, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 5, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 5, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 5, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 5, 7, 7, 7, 7, 7, 7, 7, 7}
};

 
 //code 0xe 
{{7, 7, 7, 7, 7, 7, 7, 1, 0, 0, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 1, 1, 1, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 1, 1, 1, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 1, 1, 1, 1, 0, 0, 1, 0, 7, 0, 0, 7, 7},
{7, 7, 7, 7, 7, 7, 0, 1, 1, 0, 1, 1, 1, 0, 4, 0, 0, 0, 7},
{7, 7, 7, 1, 7, 7, 0, 1, 1, 1, 0, 0, 0, 4, 4, 7, 7, 0, 0},
{7, 7, 7, 1, 0, 0, 0, 0, 1, 1, 4, 4, 4, 0, 0, 0, 7, 0, 0},
{7, 7, 7, 1, 1, 0, 0, 1, 1, 4, 4, 4, 4, 4, 0, 0, 0, 7, 0},
{7, 7, 7, 7, 1, 1, 1, 1, 0, 4, 4, 4, 4, 4, 0, 0, 0, 7, 7},
{7, 7, 7, 7, 7, 1, 0, 0, 4, 4, 4, 4, 4, 4, 7, 0, 0, 0, 7},
{7, 7, 7, 7, 7, 7, 0, 4, 4, 4, 4, 4, 4, 7, 7, 0, 0, 0, 7},
{7, 7, 7, 7, 7, 0, 4, 4, 4, 4, 4, 0, 0, 0, 7, 7, 7, 7, 7},
{7, 4, 4, 7, 7, 4, 0, 0, 0, 0, 0, 0, 4, 4, 4, 4, 4, 7, 7},
{4, 0, 4, 7, 4, 4, 4, 4, 4, 4, 4, 4, 5, 5, 4, 4, 4, 4, 7},
{4, 4, 5, 5, 4, 4, 4, 4, 4, 4, 4, 5, 5, 5, 5, 4, 4, 4, 7},
{5, 5, 5, 4, 4, 4, 4, 4, 4, 4, 5, 5, 5, 7, 5, 5, 4, 4, 4},
{5, 5, 5, 4, 4, 4, 4, 4, 4, 4, 5, 5, 5, 7, 4, 4, 4, 4, 4},
{7, 5, 5, 4, 4, 4, 4, 4, 4, 4, 4, 5, 5, 7, 7, 0, 4, 4, 4},
{7, 7, 5, 4, 4, 4, 4, 4, 4, 4, 4, 5, 5, 5, 4, 4, 4, 4, 7},
{7, 7, 7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 5, 5, 7, 7, 7},
{7, 7, 7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 7, 7, 7},
{7, 7, 7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 5, 4, 4, 4, 4, 7, 7},
{7, 7, 7, 5, 4, 4, 4, 4, 4, 4, 4, 5, 5, 5, 4, 4, 4, 7, 7},
{7, 7, 7, 5, 4, 4, 4, 4, 4, 4, 4, 5, 5, 5, 4, 4, 4, 7, 7},
{7, 7, 7, 5, 5, 5, 4, 4, 4, 4, 7, 7, 5, 4, 4, 7, 7, 7, 7},
{7, 7, 7, 7, 4, 5, 5, 5, 5, 7, 7, 7, 4, 4, 4, 4, 7, 7, 7},
{7, 7, 7, 7, 4, 5, 5, 5, 7, 7, 7, 7, 7, 4, 0, 4, 7, 7, 7},
{7, 7, 7, 7, 4, 5, 5, 5, 5, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 4, 4, 5, 5, 5, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 4, 5, 5, 5, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 4, 4, 4, 4, 5, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 4, 4, 0, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7}
};

 
 //code 0xf 
{{7, 7, 7, 7, 7, 7, 7, 7, 7, 1, 0, 0, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 1, 1, 1, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 1, 1, 1, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 1, 1, 1, 1, 0, 0, 1, 0, 7, 0, 0, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 0, 1, 1, 0, 1, 1, 1, 0, 4, 0, 0, 0, 7},
{7, 7, 7, 7, 7, 1, 7, 7, 0, 1, 1, 1, 0, 0, 0, 4, 4, 7, 7, 0, 0},
{7, 7, 7, 7, 7, 1, 0, 0, 0, 0, 1, 1, 4, 4, 4, 0, 0, 0, 7, 0, 0},
{7, 7, 7, 7, 7, 1, 1, 0, 0, 1, 1, 4, 4, 4, 4, 4, 0, 0, 0, 7, 0},
{7, 7, 7, 7, 7, 7, 1, 1, 1, 1, 0, 4, 4, 4, 4, 4, 0, 0, 0, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 1, 0, 0, 4, 4, 4, 4, 4, 4, 7, 0, 0, 0, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 0, 4, 4, 4, 4, 4, 4, 7, 7, 0, 0, 0, 7},
{7, 7, 7, 7, 7, 7, 7, 0, 4, 4, 4, 4, 4, 0, 0, 0, 7, 7, 7, 7, 7},
{7, 7, 7, 4, 4, 7, 7, 4, 0, 0, 0, 0, 0, 0, 4, 4, 4, 4, 4, 7, 7},
{7, 7, 4, 0, 4, 7, 4, 4, 4, 4, 4, 4, 4, 4, 5, 5, 4, 4, 4, 4, 7},
{7, 7, 4, 4, 5, 5, 4, 4, 4, 4, 4, 4, 4, 5, 5, 5, 5, 4, 4, 4, 7},
{7, 7, 5, 5, 5, 4, 4, 4, 4, 4, 4, 4, 5, 5, 5, 7, 5, 5, 4, 4, 4},
{7, 7, 5, 5, 5, 4, 4, 4, 4, 4, 4, 4, 5, 5, 5, 7, 4, 4, 4, 4, 4},
{7, 7, 7, 5, 5, 4, 4, 4, 4, 4, 4, 4, 4, 5, 5, 7, 7, 0, 4, 4, 4},
{7, 7, 7, 7, 5, 4, 4, 4, 4, 4, 4, 4, 4, 5, 5, 5, 4, 4, 4, 4, 7},
{4, 4, 7, 7, 7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 7, 7, 7, 7, 7, 7},
{0, 4, 7, 5, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 7, 4, 4, 7},
{4, 4, 4, 5, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 0, 7},
{0, 4, 5, 5, 5, 5, 4, 4, 4, 4, 4, 4, 4, 5, 5, 4, 4, 4, 4, 4, 7},
{7, 5, 5, 7, 5, 5, 5, 4, 4, 4, 4, 5, 5, 7, 5, 5, 5, 4, 4, 0, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 5, 4, 4, 7, 7}
};

 
 //code 0x10 
{{7, 7, 7, 7, 7, 7, 7, 1, 0, 0, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 1, 1, 1, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 1, 1, 1, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 1, 1, 1, 1, 0, 0, 1, 0, 7, 0, 0, 7, 7},
{7, 7, 7, 7, 7, 7, 0, 1, 1, 0, 1, 1, 1, 0, 4, 0, 0, 0, 7},
{7, 7, 7, 1, 7, 7, 0, 1, 1, 1, 0, 0, 0, 4, 4, 7, 7, 0, 0},
{7, 7, 7, 1, 0, 0, 0, 0, 1, 1, 4, 4, 4, 0, 0, 0, 7, 0, 0},
{7, 7, 7, 1, 1, 0, 0, 1, 1, 4, 4, 4, 4, 4, 0, 0, 0, 7, 0},
{7, 7, 7, 7, 1, 1, 1, 1, 0, 4, 4, 4, 4, 4, 0, 0, 0, 7, 7},
{7, 7, 7, 7, 7, 1, 0, 0, 4, 4, 4, 4, 4, 4, 7, 0, 0, 0, 7},
{7, 7, 7, 7, 7, 7, 0, 4, 4, 4, 4, 4, 4, 7, 7, 0, 0, 0, 7},
{7, 7, 7, 7, 7, 0, 4, 4, 4, 4, 4, 0, 0, 0, 7, 7, 7, 7, 7},
{7, 4, 4, 7, 7, 4, 0, 0, 0, 0, 0, 0, 4, 4, 4, 4, 4, 7, 7},
{4, 0, 4, 7, 4, 4, 4, 4, 4, 4, 4, 4, 5, 5, 4, 4, 4, 4, 7},
{4, 4, 5, 5, 4, 4, 4, 4, 4, 4, 4, 5, 5, 5, 5, 4, 4, 4, 7},
{5, 5, 5, 4, 4, 4, 4, 4, 4, 4, 5, 5, 5, 7, 5, 5, 4, 4, 4},
{5, 5, 5, 4, 4, 4, 4, 4, 4, 4, 5, 5, 5, 7, 4, 4, 4, 4, 4},
{7, 5, 5, 4, 4, 4, 4, 4, 4, 4, 4, 5, 5, 7, 7, 0, 4, 4, 4},
{7, 7, 5, 4, 4, 4, 4, 4, 4, 4, 4, 5, 5, 5, 4, 4, 4, 4, 7},
{7, 7, 7, 4, 4, 4, 4, 4, 4, 4, 5, 5, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 4, 4, 4, 4, 4, 4, 4, 4, 5, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 5, 4, 4, 4, 4, 4, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 4, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 7, 7, 7, 7, 7, 7},
{7, 7, 4, 5, 5, 4, 4, 4, 4, 5, 4, 4, 4, 7, 7, 7, 7, 7, 7},
{7, 7, 4, 5, 5, 5, 7, 7, 7, 5, 5, 4, 4, 7, 7, 7, 7, 7, 7},
{7, 7, 4, 4, 5, 5, 7, 7, 7, 5, 5, 4, 4, 7, 7, 7, 7, 7, 7},
{7, 7, 4, 4, 5, 5, 5, 7, 5, 5, 5, 4, 4, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 4, 4, 4, 5, 7, 5, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 4, 4, 4, 7, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 4, 0, 4, 7, 4, 0, 4, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 4, 4, 7, 7, 7, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7}
};

 
 //code 0x11 
{{7, 7, 7, 7, 7, 7, 7, 7, 4, 4, 4, 4, 4, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 4, 0, 0, 4, 0, 0, 4, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 0, 0, 4, 1, 1, 4, 1, 1, 4, 0, 0, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 0, 0, 7, 4, 1, 0, 4, 0, 1, 4, 7, 0, 0, 7, 7, 7, 7},
{7, 7, 7, 7, 0, 0, 7, 4, 1, 1, 4, 1, 1, 4, 7, 0, 0, 7, 7, 7, 7},
{7, 7, 7, 0, 0, 7, 1, 1, 1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 7, 7, 7},
{7, 7, 7, 0, 0, 1, 1, 1, 1, 1, 0, 1, 1, 1, 1, 1, 0, 0, 7, 7, 7},
{7, 7, 7, 0, 0, 1, 0, 0, 0, 1, 1, 1, 0, 0, 0, 1, 0, 0, 7, 7, 7},
{7, 7, 7, 0, 0, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 1, 0, 0, 7, 7, 7},
{7, 7, 7, 0, 7, 1, 0, 1, 0, 1, 0, 1, 0, 1, 0, 1, 7, 0, 7, 7, 7},
{7, 7, 7, 7, 7, 1, 1, 0, 0, 0, 0, 0, 0, 0, 1, 1, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 1, 1, 1, 1, 1, 1, 1, 1, 1, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 0, 4, 4, 4, 4, 4, 0, 0, 0, 7, 7, 7, 7, 7},
{7, 7, 7, 4, 4, 7, 7, 4, 0, 0, 0, 0, 0, 0, 4, 4, 4, 4, 4, 7, 7},
{7, 7, 4, 0, 4, 7, 4, 4, 4, 4, 4, 4, 4, 4, 5, 5, 4, 4, 4, 4, 7},
{7, 7, 4, 4, 5, 5, 4, 4, 4, 4, 4, 4, 4, 5, 5, 5, 5, 4, 4, 4, 7},
{7, 7, 5, 5, 5, 4, 4, 4, 4, 4, 4, 4, 5, 5, 5, 7, 5, 5, 4, 4, 4},
{7, 7, 5, 5, 5, 4, 4, 4, 4, 4, 4, 4, 5, 5, 5, 7, 4, 4, 4, 4, 4},
{7, 7, 7, 5, 5, 4, 4, 4, 4, 4, 4, 4, 4, 5, 5, 7, 7, 0, 4, 4, 4},
{7, 7, 7, 7, 5, 4, 4, 4, 4, 4, 4, 4, 4, 5, 5, 5, 4, 4, 4, 4, 7},
{4, 4, 7, 7, 7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 7, 7, 7, 7, 7, 7},
{0, 4, 7, 5, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 7, 4, 4, 7},
{4, 4, 4, 5, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 0, 7},
{0, 4, 5, 5, 5, 5, 4, 4, 4, 4, 4, 4, 4, 5, 5, 4, 4, 4, 4, 4, 7},
{7, 5, 5, 7, 5, 5, 5, 4, 4, 4, 4, 5, 5, 7, 5, 5, 5, 4, 4, 0, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 5, 4, 4, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7}
};

 
 //code 0x12 
{{7, 7, 7, 7, 0, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 0, 7, 7, 7, 7},
{7, 7, 7, 0, 0, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 0, 0, 7, 7, 7},
{7, 7, 7, 0, 0, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 0, 0, 7, 7, 7},
{7, 7, 7, 0, 0, 0, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 0, 0, 7, 7, 7},
{7, 7, 7, 0, 0, 0, 7, 7, 4, 4, 4, 4, 4, 7, 7, 0, 0, 0, 7, 7, 7},
{7, 7, 7, 7, 0, 0, 7, 4, 0, 0, 4, 0, 0, 4, 7, 0, 0, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 0, 0, 4, 1, 0, 4, 0, 1, 4, 0, 0, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 4, 1, 1, 4, 1, 1, 4, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 4, 1, 0, 0, 0, 1, 4, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 1, 1, 1, 1, 0, 1, 1, 1, 1, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 1, 1, 1, 1, 1, 0, 1, 1, 1, 1, 1, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 1, 1, 1, 1, 0, 0, 0, 1, 1, 1, 1, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 1, 1, 1, 1, 0, 0, 0, 1, 1, 1, 1, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 1, 1, 1, 1, 0, 0, 0, 1, 1, 1, 1, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 1, 1, 1, 1, 1, 1, 1, 1, 1, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 0, 4, 4, 4, 4, 4, 0, 0, 0, 7, 7, 7, 7, 7},
{7, 7, 7, 4, 4, 7, 7, 4, 0, 0, 0, 0, 0, 0, 4, 4, 4, 4, 4, 7, 7},
{7, 7, 4, 0, 4, 7, 4, 4, 4, 4, 4, 4, 4, 4, 5, 5, 4, 4, 4, 4, 7},
{7, 7, 4, 4, 5, 5, 4, 4, 4, 4, 4, 4, 4, 5, 5, 5, 5, 4, 4, 4, 7},
{7, 7, 5, 5, 5, 4, 4, 4, 4, 4, 4, 4, 5, 5, 5, 7, 5, 5, 4, 4, 4},
{7, 7, 5, 5, 5, 4, 4, 4, 4, 4, 4, 4, 5, 5, 5, 7, 4, 4, 4, 4, 4},
{7, 7, 7, 5, 5, 4, 4, 4, 4, 4, 4, 4, 4, 5, 5, 7, 7, 0, 4, 4, 4},
{7, 7, 7, 7, 5, 4, 4, 4, 4, 4, 4, 4, 4, 5, 5, 5, 4, 4, 4, 4, 7},
{4, 4, 7, 7, 7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 7, 7, 7, 7, 7, 7},
{0, 4, 7, 5, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 7, 4, 4, 7},
{4, 4, 4, 5, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 0, 7},
{0, 4, 5, 5, 5, 5, 4, 4, 4, 4, 4, 4, 4, 5, 5, 4, 4, 4, 4, 4, 7},
{7, 5, 5, 7, 5, 5, 5, 4, 4, 4, 4, 5, 5, 7, 5, 5, 5, 4, 4, 0, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 5, 4, 4, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7}
};

 
 //code 0x13 
{{7, 7, 7, 7, 7, 7, 7, 4, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 0, 0, 7, 7, 7, 7, 4, 7, 7, 4, 7, 7, 0, 0, 7, 7, 7, 7},
{7, 7, 7, 0, 0, 0, 7, 7, 4, 4, 4, 4, 7, 7, 0, 0, 0, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 0, 0, 0, 4, 0, 4, 0, 4, 0, 0, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 4, 7, 7, 7, 7, 0, 0, 0, 1, 1, 4, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 4, 7, 4, 1, 1, 0, 1, 1, 4, 7, 4, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 4, 4, 1, 0, 0, 0, 1, 4, 4, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 4, 4, 0, 0, 1, 1, 0, 1, 1, 4, 7, 7, 4, 7, 7, 7, 7},
{7, 7, 7, 4, 7, 7, 4, 0, 0, 0, 0, 0, 4, 4, 4, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 4, 0, 0, 0, 0, 0, 0, 0, 0, 4, 4, 4, 7, 7, 7, 7},
{7, 7, 7, 7, 4, 4, 4, 0, 0, 0, 1, 0, 0, 0, 0, 4, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 4, 4, 0, 0, 1, 1, 1, 0, 0, 4, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 4, 0, 0, 0, 0, 1, 0, 0, 0, 4, 4, 7, 7, 7, 7, 7},
{7, 7, 7, 4, 7, 7, 4, 0, 0, 0, 0, 0, 0, 4, 4, 7, 4, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 4, 0, 0, 4, 0, 4, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 7, 0, 4, 4, 4, 4, 4, 0, 0, 0, 7, 7, 7, 7, 7},
{7, 7, 7, 4, 4, 7, 7, 4, 0, 0, 0, 0, 0, 0, 4, 4, 4, 4, 4, 7, 7},
{7, 7, 4, 0, 4, 7, 4, 4, 4, 4, 4, 4, 4, 4, 5, 5, 4, 4, 4, 4, 7},
{7, 7, 4, 4, 5, 5, 4, 4, 4, 4, 4, 4, 4, 5, 5, 5, 5, 4, 4, 4, 7},
{7, 7, 5, 5, 5, 4, 4, 4, 4, 4, 4, 4, 5, 5, 5, 7, 5, 5, 4, 4, 4},
{7, 7, 5, 5, 5, 4, 4, 4, 4, 4, 4, 4, 5, 5, 5, 7, 4, 4, 4, 4, 4},
{7, 7, 7, 5, 5, 4, 4, 4, 4, 4, 4, 4, 4, 5, 5, 7, 7, 0, 4, 4, 4},
{7, 7, 7, 7, 5, 4, 4, 4, 4, 4, 4, 4, 4, 5, 5, 5, 4, 4, 4, 4, 7},
{4, 4, 7, 7, 7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 7, 7, 7, 7, 7, 7},
{0, 4, 7, 5, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 7, 4, 4, 7},
{4, 4, 4, 5, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 0, 7},
{0, 4, 5, 5, 5, 5, 4, 4, 4, 4, 4, 4, 4, 5, 5, 4, 4, 4, 4, 4, 7},
{7, 5, 5, 7, 5, 5, 5, 4, 4, 4, 4, 5, 5, 7, 5, 5, 5, 4, 4, 0, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 5, 4, 4, 7, 7}
};

 
 //code 0x14 
{{7, 7, 0, 0, 0, 7, 7, 4, 7, 7, 7, 0, 7, 7, 4, 7, 0, 0, 7, 7, 7},
{7, 7, 0, 0, 0, 0, 7, 7, 7, 4, 7, 0, 7, 7, 7, 0, 0, 0, 7, 7, 7},
{7, 7, 7, 7, 0, 0, 7, 7, 0, 7, 7, 0, 7, 7, 7, 0, 7, 7, 7, 7, 7},
{7, 7, 4, 7, 7, 0, 0, 7, 0, 0, 7, 0, 0, 7, 0, 0, 7, 7, 7, 7, 7},
{7, 7, 4, 7, 7, 7, 0, 0, 1, 0, 0, 0, 1, 1, 0, 7, 7, 0, 7, 7, 7},
{7, 7, 7, 7, 0, 7, 7, 1, 1, 1, 0, 1, 1, 1, 7, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 0, 1, 1, 1, 1, 0, 1, 1, 1, 1, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 4, 7, 1, 1, 1, 0, 0, 0, 1, 1, 1, 7, 4, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 0, 0, 1, 1, 1, 0, 1, 1, 1, 0, 7, 7, 4, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 0, 0, 1, 0, 0, 0, 1, 0, 0, 0, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 7, 7, 7, 7, 7, 7},
{7, 7, 7, 4, 7, 7, 0, 1, 1, 1, 1, 1, 1, 1, 0, 7, 7, 0, 7, 7, 7},
{7, 7, 7, 7, 0, 0, 1, 1, 1, 0, 1, 0, 1, 1, 1, 0, 7, 7, 7, 7, 7},
{7, 7, 4, 7, 7, 0, 1, 0, 1, 0, 1, 0, 1, 0, 1, 0, 0, 7, 7, 7, 7},
{7, 7, 4, 4, 7, 0, 1, 0, 1, 1, 1, 1, 1, 0, 1, 0, 7, 7, 7, 7, 7},
{7, 7, 7, 4, 7, 0, 1, 1, 0, 0, 0, 0, 0, 1, 1, 0, 7, 7, 7, 7, 7},
{7, 7, 7, 7, 7, 7, 0, 0, 0, 4, 0, 4, 0, 0, 0, 0, 7, 7, 7, 7, 7},
{7, 7, 7, 4, 4, 7, 7, 0, 0, 0, 0, 0, 0, 0, 4, 4, 4, 4, 4, 7, 7},
{7, 7, 4, 0, 4, 4, 4, 4, 4, 4, 4, 0, 4, 4, 5, 5, 4, 4, 4, 4, 7},
{7, 7, 4, 4, 5, 5, 4, 4, 4, 4, 4, 4, 4, 5, 5, 4, 5, 4, 4, 4, 7},
{7, 7, 5, 5, 5, 4, 4, 4, 4, 4, 4, 4, 5, 5, 5, 7, 5, 5, 4, 4, 4},
{7, 7, 5, 5, 5, 4, 4, 4, 4, 4, 4, 4, 5, 5, 5, 7, 4, 4, 4, 4, 4},
{7, 7, 7, 5, 5, 4, 4, 4, 4, 4, 4, 4, 4, 5, 5, 7, 7, 0, 4, 4, 4},
{7, 7, 7, 7, 5, 4, 4, 4, 4, 4, 4, 4, 4, 5, 5, 5, 4, 4, 4, 4, 7},
{4, 4, 7, 7, 7, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 7, 7, 7, 7, 7, 7},
{0, 4, 7, 5, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 7, 4, 4, 7},
{4, 4, 4, 5, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 0, 7},
{0, 4, 5, 5, 5, 5, 4, 4, 4, 4, 4, 4, 4, 5, 5, 4, 4, 4, 4, 4, 7},
{7, 5, 5, 7, 5, 5, 5, 4, 4, 4, 4, 5, 5, 7, 5, 5, 5, 4, 4, 0, 7},
{7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 5, 4, 4, 7, 7}
};

 
 //code 0x15 
 
 
	assign data = ROM[addr]; 
 
 endmodule  