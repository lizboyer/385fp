-- finalproject.vhd

-- Generated using ACDS version 18.1 625

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity finalproject is
	port (
		clk_clk                        : in    std_logic                     := '0';             --                     clk.clk
		hex_digits_export              : out   std_logic_vector(15 downto 0);                    --              hex_digits.export
		key_external_connection_export : in    std_logic_vector(1 downto 0)  := (others => '0'); -- key_external_connection.export
		keycode_export                 : out   std_logic_vector(7 downto 0);                     --                 keycode.export
		leds_export                    : out   std_logic_vector(13 downto 0);                    --                    leds.export
		reset_reset_n                  : in    std_logic                     := '0';             --                   reset.reset_n
		sdram_wire_addr                : out   std_logic_vector(12 downto 0);                    --              sdram_wire.addr
		sdram_wire_ba                  : out   std_logic_vector(1 downto 0);                     --                        .ba
		sdram_wire_cas_n               : out   std_logic;                                        --                        .cas_n
		sdram_wire_cke                 : out   std_logic;                                        --                        .cke
		sdram_wire_cs_n                : out   std_logic;                                        --                        .cs_n
		sdram_wire_dq                  : inout std_logic_vector(15 downto 0) := (others => '0'); --                        .dq
		sdram_wire_dqm                 : out   std_logic_vector(1 downto 0);                     --                        .dqm
		sdram_wire_ras_n               : out   std_logic;                                        --                        .ras_n
		sdram_wire_we_n                : out   std_logic;                                        --                        .we_n
		spi0_MISO                      : in    std_logic                     := '0';             --                    spi0.MISO
		spi0_MOSI                      : out   std_logic;                                        --                        .MOSI
		spi0_SCLK                      : out   std_logic;                                        --                        .SCLK
		spi0_SS_n                      : out   std_logic;                                        --                        .SS_n
		usb_gpx_export                 : in    std_logic                     := '0';             --                 usb_gpx.export
		usb_irq_export                 : in    std_logic                     := '0';             --                 usb_irq.export
		usb_rst_export                 : out   std_logic;                                        --                 usb_rst.export
		vga_port_blue                  : out   std_logic_vector(3 downto 0);                     --                vga_port.blue
		vga_port_red                   : out   std_logic_vector(3 downto 0);                     --                        .red
		vga_port_green                 : out   std_logic_vector(3 downto 0);                     --                        .green
		vga_port_hs                    : out   std_logic;                                        --                        .hs
		vga_port_vs                    : out   std_logic                                         --                        .vs
	);
end entity finalproject;

architecture rtl of finalproject is
	component finalproject_VGA_text_mode_controller_0 is
		port (
			CLK           : in  std_logic                     := 'X';             -- clk
			RESET         : in  std_logic                     := 'X';             -- reset
			AVL_ADDR      : in  std_logic_vector(9 downto 0)  := (others => 'X'); -- address
			AVL_BYTE_EN   : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			AVL_READ      : in  std_logic                     := 'X';             -- read
			AVL_READDATA  : out std_logic_vector(31 downto 0);                    -- readdata
			AVL_WRITE     : in  std_logic                     := 'X';             -- write
			AVL_WRITEDATA : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			AVL_CS        : in  std_logic                     := 'X';             -- chipselect
			blue          : out std_logic_vector(3 downto 0);                     -- blue
			red           : out std_logic_vector(3 downto 0);                     -- red
			green         : out std_logic_vector(3 downto 0);                     -- green
			hs            : out std_logic;                                        -- hs
			vs            : out std_logic                                         -- vs
		);
	end component finalproject_VGA_text_mode_controller_0;

	component finalproject_hex_digits_pio is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(15 downto 0)                     -- export
		);
	end component finalproject_hex_digits_pio;

	component finalproject_jtag_uart_0 is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component finalproject_jtag_uart_0;

	component finalproject_key is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic_vector(1 downto 0)  := (others => 'X')  -- export
		);
	end component finalproject_key;

	component finalproject_keycode is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(7 downto 0)                      -- export
		);
	end component finalproject_keycode;

	component finalproject_leds_pio is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic_vector(13 downto 0)                     -- export
		);
	end component finalproject_leds_pio;

	component finalproject_nios2_gen2_0 is
		port (
			clk                                 : in  std_logic                     := 'X';             -- clk
			reset_n                             : in  std_logic                     := 'X';             -- reset_n
			reset_req                           : in  std_logic                     := 'X';             -- reset_req
			d_address                           : out std_logic_vector(27 downto 0);                    -- address
			d_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                              : out std_logic;                                        -- read
			d_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			d_write                             : out std_logic;                                        -- write
			d_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			debug_mem_slave_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                           : out std_logic_vector(27 downto 0);                    -- address
			i_read                              : out std_logic;                                        -- read
			i_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			debug_reset_request                 : out std_logic;                                        -- reset
			debug_mem_slave_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			debug_mem_slave_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			debug_mem_slave_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			debug_mem_slave_read                : in  std_logic                     := 'X';             -- read
			debug_mem_slave_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			debug_mem_slave_waitrequest         : out std_logic;                                        -- waitrequest
			debug_mem_slave_write               : in  std_logic                     := 'X';             -- write
			debug_mem_slave_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dummy_ci_port                       : out std_logic                                         -- readra
		);
	end component finalproject_nios2_gen2_0;

	component finalproject_sdram is
		port (
			clk            : in    std_logic                     := 'X';             -- clk
			reset_n        : in    std_logic                     := 'X';             -- reset_n
			az_addr        : in    std_logic_vector(24 downto 0) := (others => 'X'); -- address
			az_be_n        : in    std_logic_vector(1 downto 0)  := (others => 'X'); -- byteenable_n
			az_cs          : in    std_logic                     := 'X';             -- chipselect
			az_data        : in    std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			az_rd_n        : in    std_logic                     := 'X';             -- read_n
			az_wr_n        : in    std_logic                     := 'X';             -- write_n
			za_data        : out   std_logic_vector(15 downto 0);                    -- readdata
			za_valid       : out   std_logic;                                        -- readdatavalid
			za_waitrequest : out   std_logic;                                        -- waitrequest
			zs_addr        : out   std_logic_vector(12 downto 0);                    -- export
			zs_ba          : out   std_logic_vector(1 downto 0);                     -- export
			zs_cas_n       : out   std_logic;                                        -- export
			zs_cke         : out   std_logic;                                        -- export
			zs_cs_n        : out   std_logic;                                        -- export
			zs_dq          : inout std_logic_vector(15 downto 0) := (others => 'X'); -- export
			zs_dqm         : out   std_logic_vector(1 downto 0);                     -- export
			zs_ras_n       : out   std_logic;                                        -- export
			zs_we_n        : out   std_logic                                         -- export
		);
	end component finalproject_sdram;

	component finalproject_sdram_pll is
		port (
			clk       : in  std_logic                     := 'X';             -- clk
			reset     : in  std_logic                     := 'X';             -- reset
			read      : in  std_logic                     := 'X';             -- read
			write     : in  std_logic                     := 'X';             -- write
			address   : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata  : out std_logic_vector(31 downto 0);                    -- readdata
			writedata : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			c0        : out std_logic;                                        -- clk
			c1        : out std_logic                                         -- clk
		);
	end component finalproject_sdram_pll;

	component finalproject_spi_0 is
		port (
			clk           : in  std_logic                     := 'X';             -- clk
			reset_n       : in  std_logic                     := 'X';             -- reset_n
			data_from_cpu : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			data_to_cpu   : out std_logic_vector(15 downto 0);                    -- readdata
			mem_addr      : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- address
			read_n        : in  std_logic                     := 'X';             -- read_n
			spi_select    : in  std_logic                     := 'X';             -- chipselect
			write_n       : in  std_logic                     := 'X';             -- write_n
			irq           : out std_logic;                                        -- irq
			MISO          : in  std_logic                     := 'X';             -- export
			MOSI          : out std_logic;                                        -- export
			SCLK          : out std_logic;                                        -- export
			SS_n          : out std_logic                                         -- export
		);
	end component finalproject_spi_0;

	component finalproject_sysid_qsys_0 is
		port (
			clock    : in  std_logic                     := 'X'; -- clk
			reset_n  : in  std_logic                     := 'X'; -- reset_n
			readdata : out std_logic_vector(31 downto 0);        -- readdata
			address  : in  std_logic                     := 'X'  -- address
		);
	end component finalproject_sysid_qsys_0;

	component finalproject_timer_0 is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- address
			writedata  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- writedata
			readdata   : out std_logic_vector(15 downto 0);                    -- readdata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write_n    : in  std_logic                     := 'X';             -- write_n
			irq        : out std_logic                                         -- irq
		);
	end component finalproject_timer_0;

	component finalproject_usb_gpx is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic                     := 'X'              -- export
		);
	end component finalproject_usb_gpx;

	component finalproject_usb_rst is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic                                         -- export
		);
	end component finalproject_usb_rst;

	component finalproject_mm_interconnect_0 is
		port (
			clk_0_clk_clk                                         : in  std_logic                     := 'X';             -- clk
			sdram_pll_c0_clk                                      : in  std_logic                     := 'X';             -- clk
			nios2_gen2_0_reset_reset_bridge_in_reset_reset        : in  std_logic                     := 'X';             -- reset
			sdram_reset_reset_bridge_in_reset_reset               : in  std_logic                     := 'X';             -- reset
			nios2_gen2_0_data_master_address                      : in  std_logic_vector(27 downto 0) := (others => 'X'); -- address
			nios2_gen2_0_data_master_waitrequest                  : out std_logic;                                        -- waitrequest
			nios2_gen2_0_data_master_byteenable                   : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			nios2_gen2_0_data_master_read                         : in  std_logic                     := 'X';             -- read
			nios2_gen2_0_data_master_readdata                     : out std_logic_vector(31 downto 0);                    -- readdata
			nios2_gen2_0_data_master_write                        : in  std_logic                     := 'X';             -- write
			nios2_gen2_0_data_master_writedata                    : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			nios2_gen2_0_data_master_debugaccess                  : in  std_logic                     := 'X';             -- debugaccess
			nios2_gen2_0_instruction_master_address               : in  std_logic_vector(27 downto 0) := (others => 'X'); -- address
			nios2_gen2_0_instruction_master_waitrequest           : out std_logic;                                        -- waitrequest
			nios2_gen2_0_instruction_master_read                  : in  std_logic                     := 'X';             -- read
			nios2_gen2_0_instruction_master_readdata              : out std_logic_vector(31 downto 0);                    -- readdata
			hex_digits_pio_s1_address                             : out std_logic_vector(1 downto 0);                     -- address
			hex_digits_pio_s1_write                               : out std_logic;                                        -- write
			hex_digits_pio_s1_readdata                            : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			hex_digits_pio_s1_writedata                           : out std_logic_vector(31 downto 0);                    -- writedata
			hex_digits_pio_s1_chipselect                          : out std_logic;                                        -- chipselect
			jtag_uart_0_avalon_jtag_slave_address                 : out std_logic_vector(0 downto 0);                     -- address
			jtag_uart_0_avalon_jtag_slave_write                   : out std_logic;                                        -- write
			jtag_uart_0_avalon_jtag_slave_read                    : out std_logic;                                        -- read
			jtag_uart_0_avalon_jtag_slave_readdata                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			jtag_uart_0_avalon_jtag_slave_writedata               : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_uart_0_avalon_jtag_slave_waitrequest             : in  std_logic                     := 'X';             -- waitrequest
			jtag_uart_0_avalon_jtag_slave_chipselect              : out std_logic;                                        -- chipselect
			key_s1_address                                        : out std_logic_vector(1 downto 0);                     -- address
			key_s1_readdata                                       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			keycode_s1_address                                    : out std_logic_vector(1 downto 0);                     -- address
			keycode_s1_write                                      : out std_logic;                                        -- write
			keycode_s1_readdata                                   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			keycode_s1_writedata                                  : out std_logic_vector(31 downto 0);                    -- writedata
			keycode_s1_chipselect                                 : out std_logic;                                        -- chipselect
			leds_pio_s1_address                                   : out std_logic_vector(1 downto 0);                     -- address
			leds_pio_s1_write                                     : out std_logic;                                        -- write
			leds_pio_s1_readdata                                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			leds_pio_s1_writedata                                 : out std_logic_vector(31 downto 0);                    -- writedata
			leds_pio_s1_chipselect                                : out std_logic;                                        -- chipselect
			nios2_gen2_0_debug_mem_slave_address                  : out std_logic_vector(8 downto 0);                     -- address
			nios2_gen2_0_debug_mem_slave_write                    : out std_logic;                                        -- write
			nios2_gen2_0_debug_mem_slave_read                     : out std_logic;                                        -- read
			nios2_gen2_0_debug_mem_slave_readdata                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			nios2_gen2_0_debug_mem_slave_writedata                : out std_logic_vector(31 downto 0);                    -- writedata
			nios2_gen2_0_debug_mem_slave_byteenable               : out std_logic_vector(3 downto 0);                     -- byteenable
			nios2_gen2_0_debug_mem_slave_waitrequest              : in  std_logic                     := 'X';             -- waitrequest
			nios2_gen2_0_debug_mem_slave_debugaccess              : out std_logic;                                        -- debugaccess
			sdram_s1_address                                      : out std_logic_vector(24 downto 0);                    -- address
			sdram_s1_write                                        : out std_logic;                                        -- write
			sdram_s1_read                                         : out std_logic;                                        -- read
			sdram_s1_readdata                                     : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			sdram_s1_writedata                                    : out std_logic_vector(15 downto 0);                    -- writedata
			sdram_s1_byteenable                                   : out std_logic_vector(1 downto 0);                     -- byteenable
			sdram_s1_readdatavalid                                : in  std_logic                     := 'X';             -- readdatavalid
			sdram_s1_waitrequest                                  : in  std_logic                     := 'X';             -- waitrequest
			sdram_s1_chipselect                                   : out std_logic;                                        -- chipselect
			sdram_pll_pll_slave_address                           : out std_logic_vector(1 downto 0);                     -- address
			sdram_pll_pll_slave_write                             : out std_logic;                                        -- write
			sdram_pll_pll_slave_read                              : out std_logic;                                        -- read
			sdram_pll_pll_slave_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			sdram_pll_pll_slave_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			spi_0_spi_control_port_address                        : out std_logic_vector(2 downto 0);                     -- address
			spi_0_spi_control_port_write                          : out std_logic;                                        -- write
			spi_0_spi_control_port_read                           : out std_logic;                                        -- read
			spi_0_spi_control_port_readdata                       : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			spi_0_spi_control_port_writedata                      : out std_logic_vector(15 downto 0);                    -- writedata
			spi_0_spi_control_port_chipselect                     : out std_logic;                                        -- chipselect
			sysid_qsys_0_control_slave_address                    : out std_logic_vector(0 downto 0);                     -- address
			sysid_qsys_0_control_slave_readdata                   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			timer_0_s1_address                                    : out std_logic_vector(3 downto 0);                     -- address
			timer_0_s1_write                                      : out std_logic;                                        -- write
			timer_0_s1_readdata                                   : in  std_logic_vector(15 downto 0) := (others => 'X'); -- readdata
			timer_0_s1_writedata                                  : out std_logic_vector(15 downto 0);                    -- writedata
			timer_0_s1_chipselect                                 : out std_logic;                                        -- chipselect
			usb_gpx_s1_address                                    : out std_logic_vector(1 downto 0);                     -- address
			usb_gpx_s1_readdata                                   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			usb_irq_s1_address                                    : out std_logic_vector(1 downto 0);                     -- address
			usb_irq_s1_readdata                                   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			usb_rst_s1_address                                    : out std_logic_vector(1 downto 0);                     -- address
			usb_rst_s1_write                                      : out std_logic;                                        -- write
			usb_rst_s1_readdata                                   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			usb_rst_s1_writedata                                  : out std_logic_vector(31 downto 0);                    -- writedata
			usb_rst_s1_chipselect                                 : out std_logic;                                        -- chipselect
			VGA_text_mode_controller_0_avalon_mm_slave_address    : out std_logic_vector(9 downto 0);                     -- address
			VGA_text_mode_controller_0_avalon_mm_slave_write      : out std_logic;                                        -- write
			VGA_text_mode_controller_0_avalon_mm_slave_read       : out std_logic;                                        -- read
			VGA_text_mode_controller_0_avalon_mm_slave_readdata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			VGA_text_mode_controller_0_avalon_mm_slave_writedata  : out std_logic_vector(31 downto 0);                    -- writedata
			VGA_text_mode_controller_0_avalon_mm_slave_byteenable : out std_logic_vector(3 downto 0);                     -- byteenable
			VGA_text_mode_controller_0_avalon_mm_slave_chipselect : out std_logic                                         -- chipselect
		);
	end component finalproject_mm_interconnect_0;

	component finalproject_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			receiver1_irq : in  std_logic                     := 'X'; -- irq
			receiver2_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component finalproject_irq_mapper;

	component finalproject_rst_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			reset_in1      : in  std_logic := 'X'; -- reset_in1.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_req      : out std_logic;        --          .reset_req
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component finalproject_rst_controller;

	component finalproject_rst_controller_001 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			reset_in1      : in  std_logic := 'X'; -- reset_in1.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req      : out std_logic;
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component finalproject_rst_controller_001;

	signal sdram_pll_c0_clk                                                        : std_logic;                     -- sdram_pll:c0 -> [mm_interconnect_0:sdram_pll_c0_clk, rst_controller_001:clk, sdram:clk]
	signal nios2_gen2_0_data_master_readdata                                       : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_gen2_0_data_master_readdata -> nios2_gen2_0:d_readdata
	signal nios2_gen2_0_data_master_waitrequest                                    : std_logic;                     -- mm_interconnect_0:nios2_gen2_0_data_master_waitrequest -> nios2_gen2_0:d_waitrequest
	signal nios2_gen2_0_data_master_debugaccess                                    : std_logic;                     -- nios2_gen2_0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_gen2_0_data_master_debugaccess
	signal nios2_gen2_0_data_master_address                                        : std_logic_vector(27 downto 0); -- nios2_gen2_0:d_address -> mm_interconnect_0:nios2_gen2_0_data_master_address
	signal nios2_gen2_0_data_master_byteenable                                     : std_logic_vector(3 downto 0);  -- nios2_gen2_0:d_byteenable -> mm_interconnect_0:nios2_gen2_0_data_master_byteenable
	signal nios2_gen2_0_data_master_read                                           : std_logic;                     -- nios2_gen2_0:d_read -> mm_interconnect_0:nios2_gen2_0_data_master_read
	signal nios2_gen2_0_data_master_write                                          : std_logic;                     -- nios2_gen2_0:d_write -> mm_interconnect_0:nios2_gen2_0_data_master_write
	signal nios2_gen2_0_data_master_writedata                                      : std_logic_vector(31 downto 0); -- nios2_gen2_0:d_writedata -> mm_interconnect_0:nios2_gen2_0_data_master_writedata
	signal nios2_gen2_0_instruction_master_readdata                                : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_gen2_0_instruction_master_readdata -> nios2_gen2_0:i_readdata
	signal nios2_gen2_0_instruction_master_waitrequest                             : std_logic;                     -- mm_interconnect_0:nios2_gen2_0_instruction_master_waitrequest -> nios2_gen2_0:i_waitrequest
	signal nios2_gen2_0_instruction_master_address                                 : std_logic_vector(27 downto 0); -- nios2_gen2_0:i_address -> mm_interconnect_0:nios2_gen2_0_instruction_master_address
	signal nios2_gen2_0_instruction_master_read                                    : std_logic;                     -- nios2_gen2_0:i_read -> mm_interconnect_0:nios2_gen2_0_instruction_master_read
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect              : std_logic;                     -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata                : std_logic_vector(31 downto 0); -- jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest             : std_logic;                     -- jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address                 : std_logic_vector(0 downto 0);  -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read                    : std_logic;                     -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read:in
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write                   : std_logic;                     -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write:in
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata               : std_logic_vector(31 downto 0); -- mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	signal mm_interconnect_0_vga_text_mode_controller_0_avalon_mm_slave_chipselect : std_logic;                     -- mm_interconnect_0:VGA_text_mode_controller_0_avalon_mm_slave_chipselect -> VGA_text_mode_controller_0:AVL_CS
	signal mm_interconnect_0_vga_text_mode_controller_0_avalon_mm_slave_readdata   : std_logic_vector(31 downto 0); -- VGA_text_mode_controller_0:AVL_READDATA -> mm_interconnect_0:VGA_text_mode_controller_0_avalon_mm_slave_readdata
	signal mm_interconnect_0_vga_text_mode_controller_0_avalon_mm_slave_address    : std_logic_vector(9 downto 0);  -- mm_interconnect_0:VGA_text_mode_controller_0_avalon_mm_slave_address -> VGA_text_mode_controller_0:AVL_ADDR
	signal mm_interconnect_0_vga_text_mode_controller_0_avalon_mm_slave_read       : std_logic;                     -- mm_interconnect_0:VGA_text_mode_controller_0_avalon_mm_slave_read -> VGA_text_mode_controller_0:AVL_READ
	signal mm_interconnect_0_vga_text_mode_controller_0_avalon_mm_slave_byteenable : std_logic_vector(3 downto 0);  -- mm_interconnect_0:VGA_text_mode_controller_0_avalon_mm_slave_byteenable -> VGA_text_mode_controller_0:AVL_BYTE_EN
	signal mm_interconnect_0_vga_text_mode_controller_0_avalon_mm_slave_write      : std_logic;                     -- mm_interconnect_0:VGA_text_mode_controller_0_avalon_mm_slave_write -> VGA_text_mode_controller_0:AVL_WRITE
	signal mm_interconnect_0_vga_text_mode_controller_0_avalon_mm_slave_writedata  : std_logic_vector(31 downto 0); -- mm_interconnect_0:VGA_text_mode_controller_0_avalon_mm_slave_writedata -> VGA_text_mode_controller_0:AVL_WRITEDATA
	signal mm_interconnect_0_sysid_qsys_0_control_slave_readdata                   : std_logic_vector(31 downto 0); -- sysid_qsys_0:readdata -> mm_interconnect_0:sysid_qsys_0_control_slave_readdata
	signal mm_interconnect_0_sysid_qsys_0_control_slave_address                    : std_logic_vector(0 downto 0);  -- mm_interconnect_0:sysid_qsys_0_control_slave_address -> sysid_qsys_0:address
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata                 : std_logic_vector(31 downto 0); -- nios2_gen2_0:debug_mem_slave_readdata -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_readdata
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest              : std_logic;                     -- nios2_gen2_0:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_waitrequest
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess              : std_logic;                     -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_debugaccess -> nios2_gen2_0:debug_mem_slave_debugaccess
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address                  : std_logic_vector(8 downto 0);  -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_address -> nios2_gen2_0:debug_mem_slave_address
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read                     : std_logic;                     -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_read -> nios2_gen2_0:debug_mem_slave_read
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable               : std_logic_vector(3 downto 0);  -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_byteenable -> nios2_gen2_0:debug_mem_slave_byteenable
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write                    : std_logic;                     -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_write -> nios2_gen2_0:debug_mem_slave_write
	signal mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata                : std_logic_vector(31 downto 0); -- mm_interconnect_0:nios2_gen2_0_debug_mem_slave_writedata -> nios2_gen2_0:debug_mem_slave_writedata
	signal mm_interconnect_0_sdram_pll_pll_slave_readdata                          : std_logic_vector(31 downto 0); -- sdram_pll:readdata -> mm_interconnect_0:sdram_pll_pll_slave_readdata
	signal mm_interconnect_0_sdram_pll_pll_slave_address                           : std_logic_vector(1 downto 0);  -- mm_interconnect_0:sdram_pll_pll_slave_address -> sdram_pll:address
	signal mm_interconnect_0_sdram_pll_pll_slave_read                              : std_logic;                     -- mm_interconnect_0:sdram_pll_pll_slave_read -> sdram_pll:read
	signal mm_interconnect_0_sdram_pll_pll_slave_write                             : std_logic;                     -- mm_interconnect_0:sdram_pll_pll_slave_write -> sdram_pll:write
	signal mm_interconnect_0_sdram_pll_pll_slave_writedata                         : std_logic_vector(31 downto 0); -- mm_interconnect_0:sdram_pll_pll_slave_writedata -> sdram_pll:writedata
	signal mm_interconnect_0_sdram_s1_chipselect                                   : std_logic;                     -- mm_interconnect_0:sdram_s1_chipselect -> sdram:az_cs
	signal mm_interconnect_0_sdram_s1_readdata                                     : std_logic_vector(15 downto 0); -- sdram:za_data -> mm_interconnect_0:sdram_s1_readdata
	signal mm_interconnect_0_sdram_s1_waitrequest                                  : std_logic;                     -- sdram:za_waitrequest -> mm_interconnect_0:sdram_s1_waitrequest
	signal mm_interconnect_0_sdram_s1_address                                      : std_logic_vector(24 downto 0); -- mm_interconnect_0:sdram_s1_address -> sdram:az_addr
	signal mm_interconnect_0_sdram_s1_read                                         : std_logic;                     -- mm_interconnect_0:sdram_s1_read -> mm_interconnect_0_sdram_s1_read:in
	signal mm_interconnect_0_sdram_s1_byteenable                                   : std_logic_vector(1 downto 0);  -- mm_interconnect_0:sdram_s1_byteenable -> mm_interconnect_0_sdram_s1_byteenable:in
	signal mm_interconnect_0_sdram_s1_readdatavalid                                : std_logic;                     -- sdram:za_valid -> mm_interconnect_0:sdram_s1_readdatavalid
	signal mm_interconnect_0_sdram_s1_write                                        : std_logic;                     -- mm_interconnect_0:sdram_s1_write -> mm_interconnect_0_sdram_s1_write:in
	signal mm_interconnect_0_sdram_s1_writedata                                    : std_logic_vector(15 downto 0); -- mm_interconnect_0:sdram_s1_writedata -> sdram:az_data
	signal mm_interconnect_0_keycode_s1_chipselect                                 : std_logic;                     -- mm_interconnect_0:keycode_s1_chipselect -> keycode:chipselect
	signal mm_interconnect_0_keycode_s1_readdata                                   : std_logic_vector(31 downto 0); -- keycode:readdata -> mm_interconnect_0:keycode_s1_readdata
	signal mm_interconnect_0_keycode_s1_address                                    : std_logic_vector(1 downto 0);  -- mm_interconnect_0:keycode_s1_address -> keycode:address
	signal mm_interconnect_0_keycode_s1_write                                      : std_logic;                     -- mm_interconnect_0:keycode_s1_write -> mm_interconnect_0_keycode_s1_write:in
	signal mm_interconnect_0_keycode_s1_writedata                                  : std_logic_vector(31 downto 0); -- mm_interconnect_0:keycode_s1_writedata -> keycode:writedata
	signal mm_interconnect_0_usb_irq_s1_readdata                                   : std_logic_vector(31 downto 0); -- usb_irq:readdata -> mm_interconnect_0:usb_irq_s1_readdata
	signal mm_interconnect_0_usb_irq_s1_address                                    : std_logic_vector(1 downto 0);  -- mm_interconnect_0:usb_irq_s1_address -> usb_irq:address
	signal mm_interconnect_0_usb_gpx_s1_readdata                                   : std_logic_vector(31 downto 0); -- usb_gpx:readdata -> mm_interconnect_0:usb_gpx_s1_readdata
	signal mm_interconnect_0_usb_gpx_s1_address                                    : std_logic_vector(1 downto 0);  -- mm_interconnect_0:usb_gpx_s1_address -> usb_gpx:address
	signal mm_interconnect_0_usb_rst_s1_chipselect                                 : std_logic;                     -- mm_interconnect_0:usb_rst_s1_chipselect -> usb_rst:chipselect
	signal mm_interconnect_0_usb_rst_s1_readdata                                   : std_logic_vector(31 downto 0); -- usb_rst:readdata -> mm_interconnect_0:usb_rst_s1_readdata
	signal mm_interconnect_0_usb_rst_s1_address                                    : std_logic_vector(1 downto 0);  -- mm_interconnect_0:usb_rst_s1_address -> usb_rst:address
	signal mm_interconnect_0_usb_rst_s1_write                                      : std_logic;                     -- mm_interconnect_0:usb_rst_s1_write -> mm_interconnect_0_usb_rst_s1_write:in
	signal mm_interconnect_0_usb_rst_s1_writedata                                  : std_logic_vector(31 downto 0); -- mm_interconnect_0:usb_rst_s1_writedata -> usb_rst:writedata
	signal mm_interconnect_0_hex_digits_pio_s1_chipselect                          : std_logic;                     -- mm_interconnect_0:hex_digits_pio_s1_chipselect -> hex_digits_pio:chipselect
	signal mm_interconnect_0_hex_digits_pio_s1_readdata                            : std_logic_vector(31 downto 0); -- hex_digits_pio:readdata -> mm_interconnect_0:hex_digits_pio_s1_readdata
	signal mm_interconnect_0_hex_digits_pio_s1_address                             : std_logic_vector(1 downto 0);  -- mm_interconnect_0:hex_digits_pio_s1_address -> hex_digits_pio:address
	signal mm_interconnect_0_hex_digits_pio_s1_write                               : std_logic;                     -- mm_interconnect_0:hex_digits_pio_s1_write -> mm_interconnect_0_hex_digits_pio_s1_write:in
	signal mm_interconnect_0_hex_digits_pio_s1_writedata                           : std_logic_vector(31 downto 0); -- mm_interconnect_0:hex_digits_pio_s1_writedata -> hex_digits_pio:writedata
	signal mm_interconnect_0_leds_pio_s1_chipselect                                : std_logic;                     -- mm_interconnect_0:leds_pio_s1_chipselect -> leds_pio:chipselect
	signal mm_interconnect_0_leds_pio_s1_readdata                                  : std_logic_vector(31 downto 0); -- leds_pio:readdata -> mm_interconnect_0:leds_pio_s1_readdata
	signal mm_interconnect_0_leds_pio_s1_address                                   : std_logic_vector(1 downto 0);  -- mm_interconnect_0:leds_pio_s1_address -> leds_pio:address
	signal mm_interconnect_0_leds_pio_s1_write                                     : std_logic;                     -- mm_interconnect_0:leds_pio_s1_write -> mm_interconnect_0_leds_pio_s1_write:in
	signal mm_interconnect_0_leds_pio_s1_writedata                                 : std_logic_vector(31 downto 0); -- mm_interconnect_0:leds_pio_s1_writedata -> leds_pio:writedata
	signal mm_interconnect_0_key_s1_readdata                                       : std_logic_vector(31 downto 0); -- key:readdata -> mm_interconnect_0:key_s1_readdata
	signal mm_interconnect_0_key_s1_address                                        : std_logic_vector(1 downto 0);  -- mm_interconnect_0:key_s1_address -> key:address
	signal mm_interconnect_0_timer_0_s1_chipselect                                 : std_logic;                     -- mm_interconnect_0:timer_0_s1_chipselect -> timer_0:chipselect
	signal mm_interconnect_0_timer_0_s1_readdata                                   : std_logic_vector(15 downto 0); -- timer_0:readdata -> mm_interconnect_0:timer_0_s1_readdata
	signal mm_interconnect_0_timer_0_s1_address                                    : std_logic_vector(3 downto 0);  -- mm_interconnect_0:timer_0_s1_address -> timer_0:address
	signal mm_interconnect_0_timer_0_s1_write                                      : std_logic;                     -- mm_interconnect_0:timer_0_s1_write -> mm_interconnect_0_timer_0_s1_write:in
	signal mm_interconnect_0_timer_0_s1_writedata                                  : std_logic_vector(15 downto 0); -- mm_interconnect_0:timer_0_s1_writedata -> timer_0:writedata
	signal mm_interconnect_0_spi_0_spi_control_port_chipselect                     : std_logic;                     -- mm_interconnect_0:spi_0_spi_control_port_chipselect -> spi_0:spi_select
	signal mm_interconnect_0_spi_0_spi_control_port_readdata                       : std_logic_vector(15 downto 0); -- spi_0:data_to_cpu -> mm_interconnect_0:spi_0_spi_control_port_readdata
	signal mm_interconnect_0_spi_0_spi_control_port_address                        : std_logic_vector(2 downto 0);  -- mm_interconnect_0:spi_0_spi_control_port_address -> spi_0:mem_addr
	signal mm_interconnect_0_spi_0_spi_control_port_read                           : std_logic;                     -- mm_interconnect_0:spi_0_spi_control_port_read -> mm_interconnect_0_spi_0_spi_control_port_read:in
	signal mm_interconnect_0_spi_0_spi_control_port_write                          : std_logic;                     -- mm_interconnect_0:spi_0_spi_control_port_write -> mm_interconnect_0_spi_0_spi_control_port_write:in
	signal mm_interconnect_0_spi_0_spi_control_port_writedata                      : std_logic_vector(15 downto 0); -- mm_interconnect_0:spi_0_spi_control_port_writedata -> spi_0:data_from_cpu
	signal irq_mapper_receiver0_irq                                                : std_logic;                     -- jtag_uart_0:av_irq -> irq_mapper:receiver0_irq
	signal irq_mapper_receiver1_irq                                                : std_logic;                     -- timer_0:irq -> irq_mapper:receiver1_irq
	signal irq_mapper_receiver2_irq                                                : std_logic;                     -- spi_0:irq -> irq_mapper:receiver2_irq
	signal nios2_gen2_0_irq_irq                                                    : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> nios2_gen2_0:irq
	signal rst_controller_reset_out_reset                                          : std_logic;                     -- rst_controller:reset_out -> [VGA_text_mode_controller_0:RESET, irq_mapper:reset, mm_interconnect_0:nios2_gen2_0_reset_reset_bridge_in_reset_reset, rst_controller_reset_out_reset:in, rst_translator:in_reset, sdram_pll:reset]
	signal rst_controller_reset_out_reset_req                                      : std_logic;                     -- rst_controller:reset_req -> [nios2_gen2_0:reset_req, rst_translator:reset_req_in]
	signal nios2_gen2_0_debug_reset_request_reset                                  : std_logic;                     -- nios2_gen2_0:debug_reset_request -> [rst_controller:reset_in1, rst_controller_001:reset_in1]
	signal rst_controller_001_reset_out_reset                                      : std_logic;                     -- rst_controller_001:reset_out -> [mm_interconnect_0:sdram_reset_reset_bridge_in_reset_reset, rst_controller_001_reset_out_reset:in]
	signal reset_reset_n_ports_inv                                                 : std_logic;                     -- reset_reset_n:inv -> [rst_controller:reset_in0, rst_controller_001:reset_in0]
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read_ports_inv          : std_logic;                     -- mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read:inv -> jtag_uart_0:av_read_n
	signal mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write_ports_inv         : std_logic;                     -- mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write:inv -> jtag_uart_0:av_write_n
	signal mm_interconnect_0_sdram_s1_read_ports_inv                               : std_logic;                     -- mm_interconnect_0_sdram_s1_read:inv -> sdram:az_rd_n
	signal mm_interconnect_0_sdram_s1_byteenable_ports_inv                         : std_logic_vector(1 downto 0);  -- mm_interconnect_0_sdram_s1_byteenable:inv -> sdram:az_be_n
	signal mm_interconnect_0_sdram_s1_write_ports_inv                              : std_logic;                     -- mm_interconnect_0_sdram_s1_write:inv -> sdram:az_wr_n
	signal mm_interconnect_0_keycode_s1_write_ports_inv                            : std_logic;                     -- mm_interconnect_0_keycode_s1_write:inv -> keycode:write_n
	signal mm_interconnect_0_usb_rst_s1_write_ports_inv                            : std_logic;                     -- mm_interconnect_0_usb_rst_s1_write:inv -> usb_rst:write_n
	signal mm_interconnect_0_hex_digits_pio_s1_write_ports_inv                     : std_logic;                     -- mm_interconnect_0_hex_digits_pio_s1_write:inv -> hex_digits_pio:write_n
	signal mm_interconnect_0_leds_pio_s1_write_ports_inv                           : std_logic;                     -- mm_interconnect_0_leds_pio_s1_write:inv -> leds_pio:write_n
	signal mm_interconnect_0_timer_0_s1_write_ports_inv                            : std_logic;                     -- mm_interconnect_0_timer_0_s1_write:inv -> timer_0:write_n
	signal mm_interconnect_0_spi_0_spi_control_port_read_ports_inv                 : std_logic;                     -- mm_interconnect_0_spi_0_spi_control_port_read:inv -> spi_0:read_n
	signal mm_interconnect_0_spi_0_spi_control_port_write_ports_inv                : std_logic;                     -- mm_interconnect_0_spi_0_spi_control_port_write:inv -> spi_0:write_n
	signal rst_controller_reset_out_reset_ports_inv                                : std_logic;                     -- rst_controller_reset_out_reset:inv -> [hex_digits_pio:reset_n, jtag_uart_0:rst_n, key:reset_n, keycode:reset_n, leds_pio:reset_n, nios2_gen2_0:reset_n, spi_0:reset_n, sysid_qsys_0:reset_n, timer_0:reset_n, usb_gpx:reset_n, usb_irq:reset_n, usb_rst:reset_n]
	signal rst_controller_001_reset_out_reset_ports_inv                            : std_logic;                     -- rst_controller_001_reset_out_reset:inv -> sdram:reset_n

begin

	vga_text_mode_controller_0 : component finalproject_VGA_text_mode_controller_0
		port map (
			CLK           => clk_clk,                                                                 --             CLK.clk
			RESET         => rst_controller_reset_out_reset,                                          --           RESET.reset
			AVL_ADDR      => mm_interconnect_0_vga_text_mode_controller_0_avalon_mm_slave_address,    -- avalon_mm_slave.address
			AVL_BYTE_EN   => mm_interconnect_0_vga_text_mode_controller_0_avalon_mm_slave_byteenable, --                .byteenable
			AVL_READ      => mm_interconnect_0_vga_text_mode_controller_0_avalon_mm_slave_read,       --                .read
			AVL_READDATA  => mm_interconnect_0_vga_text_mode_controller_0_avalon_mm_slave_readdata,   --                .readdata
			AVL_WRITE     => mm_interconnect_0_vga_text_mode_controller_0_avalon_mm_slave_write,      --                .write
			AVL_WRITEDATA => mm_interconnect_0_vga_text_mode_controller_0_avalon_mm_slave_writedata,  --                .writedata
			AVL_CS        => mm_interconnect_0_vga_text_mode_controller_0_avalon_mm_slave_chipselect, --                .chipselect
			blue          => vga_port_blue,                                                           --        VGA_port.blue
			red           => vga_port_red,                                                            --                .red
			green         => vga_port_green,                                                          --                .green
			hs            => vga_port_hs,                                                             --                .hs
			vs            => vga_port_vs                                                              --                .vs
		);

	hex_digits_pio : component finalproject_hex_digits_pio
		port map (
			clk        => clk_clk,                                             --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,            --               reset.reset_n
			address    => mm_interconnect_0_hex_digits_pio_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_hex_digits_pio_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_hex_digits_pio_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_hex_digits_pio_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_hex_digits_pio_s1_readdata,        --                    .readdata
			out_port   => hex_digits_export                                    -- external_connection.export
		);

	jtag_uart_0 : component finalproject_jtag_uart_0
		port map (
			clk            => clk_clk,                                                         --               clk.clk
			rst_n          => rst_controller_reset_out_reset_ports_inv,                        --             reset.reset_n
			av_chipselect  => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_receiver0_irq                                         --               irq.irq
		);

	key : component finalproject_key
		port map (
			clk      => clk_clk,                                  --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv, --               reset.reset_n
			address  => mm_interconnect_0_key_s1_address,         --                  s1.address
			readdata => mm_interconnect_0_key_s1_readdata,        --                    .readdata
			in_port  => key_external_connection_export            -- external_connection.export
		);

	keycode : component finalproject_keycode
		port map (
			clk        => clk_clk,                                      --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,     --               reset.reset_n
			address    => mm_interconnect_0_keycode_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_keycode_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_keycode_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_keycode_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_keycode_s1_readdata,        --                    .readdata
			out_port   => keycode_export                                -- external_connection.export
		);

	leds_pio : component finalproject_leds_pio
		port map (
			clk        => clk_clk,                                       --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,      --               reset.reset_n
			address    => mm_interconnect_0_leds_pio_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_leds_pio_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_leds_pio_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_leds_pio_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_leds_pio_s1_readdata,        --                    .readdata
			out_port   => leds_export                                    -- external_connection.export
		);

	nios2_gen2_0 : component finalproject_nios2_gen2_0
		port map (
			clk                                 => clk_clk,                                                    --                       clk.clk
			reset_n                             => rst_controller_reset_out_reset_ports_inv,                   --                     reset.reset_n
			reset_req                           => rst_controller_reset_out_reset_req,                         --                          .reset_req
			d_address                           => nios2_gen2_0_data_master_address,                           --               data_master.address
			d_byteenable                        => nios2_gen2_0_data_master_byteenable,                        --                          .byteenable
			d_read                              => nios2_gen2_0_data_master_read,                              --                          .read
			d_readdata                          => nios2_gen2_0_data_master_readdata,                          --                          .readdata
			d_waitrequest                       => nios2_gen2_0_data_master_waitrequest,                       --                          .waitrequest
			d_write                             => nios2_gen2_0_data_master_write,                             --                          .write
			d_writedata                         => nios2_gen2_0_data_master_writedata,                         --                          .writedata
			debug_mem_slave_debugaccess_to_roms => nios2_gen2_0_data_master_debugaccess,                       --                          .debugaccess
			i_address                           => nios2_gen2_0_instruction_master_address,                    --        instruction_master.address
			i_read                              => nios2_gen2_0_instruction_master_read,                       --                          .read
			i_readdata                          => nios2_gen2_0_instruction_master_readdata,                   --                          .readdata
			i_waitrequest                       => nios2_gen2_0_instruction_master_waitrequest,                --                          .waitrequest
			irq                                 => nios2_gen2_0_irq_irq,                                       --                       irq.irq
			debug_reset_request                 => nios2_gen2_0_debug_reset_request_reset,                     --       debug_reset_request.reset
			debug_mem_slave_address             => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address,     --           debug_mem_slave.address
			debug_mem_slave_byteenable          => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable,  --                          .byteenable
			debug_mem_slave_debugaccess         => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess, --                          .debugaccess
			debug_mem_slave_read                => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read,        --                          .read
			debug_mem_slave_readdata            => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata,    --                          .readdata
			debug_mem_slave_waitrequest         => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest, --                          .waitrequest
			debug_mem_slave_write               => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write,       --                          .write
			debug_mem_slave_writedata           => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata,   --                          .writedata
			dummy_ci_port                       => open                                                        -- custom_instruction_master.readra
		);

	sdram : component finalproject_sdram
		port map (
			clk            => sdram_pll_c0_clk,                                --   clk.clk
			reset_n        => rst_controller_001_reset_out_reset_ports_inv,    -- reset.reset_n
			az_addr        => mm_interconnect_0_sdram_s1_address,              --    s1.address
			az_be_n        => mm_interconnect_0_sdram_s1_byteenable_ports_inv, --      .byteenable_n
			az_cs          => mm_interconnect_0_sdram_s1_chipselect,           --      .chipselect
			az_data        => mm_interconnect_0_sdram_s1_writedata,            --      .writedata
			az_rd_n        => mm_interconnect_0_sdram_s1_read_ports_inv,       --      .read_n
			az_wr_n        => mm_interconnect_0_sdram_s1_write_ports_inv,      --      .write_n
			za_data        => mm_interconnect_0_sdram_s1_readdata,             --      .readdata
			za_valid       => mm_interconnect_0_sdram_s1_readdatavalid,        --      .readdatavalid
			za_waitrequest => mm_interconnect_0_sdram_s1_waitrequest,          --      .waitrequest
			zs_addr        => sdram_wire_addr,                                 --  wire.export
			zs_ba          => sdram_wire_ba,                                   --      .export
			zs_cas_n       => sdram_wire_cas_n,                                --      .export
			zs_cke         => sdram_wire_cke,                                  --      .export
			zs_cs_n        => sdram_wire_cs_n,                                 --      .export
			zs_dq          => sdram_wire_dq,                                   --      .export
			zs_dqm         => sdram_wire_dqm,                                  --      .export
			zs_ras_n       => sdram_wire_ras_n,                                --      .export
			zs_we_n        => sdram_wire_we_n                                  --      .export
		);

	sdram_pll : component finalproject_sdram_pll
		port map (
			clk       => clk_clk,                                         --       inclk_interface.clk
			reset     => rst_controller_reset_out_reset,                  -- inclk_interface_reset.reset
			read      => mm_interconnect_0_sdram_pll_pll_slave_read,      --             pll_slave.read
			write     => mm_interconnect_0_sdram_pll_pll_slave_write,     --                      .write
			address   => mm_interconnect_0_sdram_pll_pll_slave_address,   --                      .address
			readdata  => mm_interconnect_0_sdram_pll_pll_slave_readdata,  --                      .readdata
			writedata => mm_interconnect_0_sdram_pll_pll_slave_writedata, --                      .writedata
			c0        => sdram_pll_c0_clk,                                --                    c0.clk
			c1        => open                                             --                    c1.clk
		);

	spi_0 : component finalproject_spi_0
		port map (
			clk           => clk_clk,                                                  --              clk.clk
			reset_n       => rst_controller_reset_out_reset_ports_inv,                 --            reset.reset_n
			data_from_cpu => mm_interconnect_0_spi_0_spi_control_port_writedata,       -- spi_control_port.writedata
			data_to_cpu   => mm_interconnect_0_spi_0_spi_control_port_readdata,        --                 .readdata
			mem_addr      => mm_interconnect_0_spi_0_spi_control_port_address,         --                 .address
			read_n        => mm_interconnect_0_spi_0_spi_control_port_read_ports_inv,  --                 .read_n
			spi_select    => mm_interconnect_0_spi_0_spi_control_port_chipselect,      --                 .chipselect
			write_n       => mm_interconnect_0_spi_0_spi_control_port_write_ports_inv, --                 .write_n
			irq           => irq_mapper_receiver2_irq,                                 --              irq.irq
			MISO          => spi0_MISO,                                                --         external.export
			MOSI          => spi0_MOSI,                                                --                 .export
			SCLK          => spi0_SCLK,                                                --                 .export
			SS_n          => spi0_SS_n                                                 --                 .export
		);

	sysid_qsys_0 : component finalproject_sysid_qsys_0
		port map (
			clock    => clk_clk,                                                 --           clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,                --         reset.reset_n
			readdata => mm_interconnect_0_sysid_qsys_0_control_slave_readdata,   -- control_slave.readdata
			address  => mm_interconnect_0_sysid_qsys_0_control_slave_address(0)  --              .address
		);

	timer_0 : component finalproject_timer_0
		port map (
			clk        => clk_clk,                                      --   clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,     -- reset.reset_n
			address    => mm_interconnect_0_timer_0_s1_address,         --    s1.address
			writedata  => mm_interconnect_0_timer_0_s1_writedata,       --      .writedata
			readdata   => mm_interconnect_0_timer_0_s1_readdata,        --      .readdata
			chipselect => mm_interconnect_0_timer_0_s1_chipselect,      --      .chipselect
			write_n    => mm_interconnect_0_timer_0_s1_write_ports_inv, --      .write_n
			irq        => irq_mapper_receiver1_irq                      --   irq.irq
		);

	usb_gpx : component finalproject_usb_gpx
		port map (
			clk      => clk_clk,                                  --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv, --               reset.reset_n
			address  => mm_interconnect_0_usb_gpx_s1_address,     --                  s1.address
			readdata => mm_interconnect_0_usb_gpx_s1_readdata,    --                    .readdata
			in_port  => usb_gpx_export                            -- external_connection.export
		);

	usb_irq : component finalproject_usb_gpx
		port map (
			clk      => clk_clk,                                  --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv, --               reset.reset_n
			address  => mm_interconnect_0_usb_irq_s1_address,     --                  s1.address
			readdata => mm_interconnect_0_usb_irq_s1_readdata,    --                    .readdata
			in_port  => usb_irq_export                            -- external_connection.export
		);

	usb_rst : component finalproject_usb_rst
		port map (
			clk        => clk_clk,                                      --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,     --               reset.reset_n
			address    => mm_interconnect_0_usb_rst_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_usb_rst_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_usb_rst_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_usb_rst_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_usb_rst_s1_readdata,        --                    .readdata
			out_port   => usb_rst_export                                -- external_connection.export
		);

	mm_interconnect_0 : component finalproject_mm_interconnect_0
		port map (
			clk_0_clk_clk                                         => clk_clk,                                                                 --                                  clk_0_clk.clk
			sdram_pll_c0_clk                                      => sdram_pll_c0_clk,                                                        --                               sdram_pll_c0.clk
			nios2_gen2_0_reset_reset_bridge_in_reset_reset        => rst_controller_reset_out_reset,                                          --   nios2_gen2_0_reset_reset_bridge_in_reset.reset
			sdram_reset_reset_bridge_in_reset_reset               => rst_controller_001_reset_out_reset,                                      --          sdram_reset_reset_bridge_in_reset.reset
			nios2_gen2_0_data_master_address                      => nios2_gen2_0_data_master_address,                                        --                   nios2_gen2_0_data_master.address
			nios2_gen2_0_data_master_waitrequest                  => nios2_gen2_0_data_master_waitrequest,                                    --                                           .waitrequest
			nios2_gen2_0_data_master_byteenable                   => nios2_gen2_0_data_master_byteenable,                                     --                                           .byteenable
			nios2_gen2_0_data_master_read                         => nios2_gen2_0_data_master_read,                                           --                                           .read
			nios2_gen2_0_data_master_readdata                     => nios2_gen2_0_data_master_readdata,                                       --                                           .readdata
			nios2_gen2_0_data_master_write                        => nios2_gen2_0_data_master_write,                                          --                                           .write
			nios2_gen2_0_data_master_writedata                    => nios2_gen2_0_data_master_writedata,                                      --                                           .writedata
			nios2_gen2_0_data_master_debugaccess                  => nios2_gen2_0_data_master_debugaccess,                                    --                                           .debugaccess
			nios2_gen2_0_instruction_master_address               => nios2_gen2_0_instruction_master_address,                                 --            nios2_gen2_0_instruction_master.address
			nios2_gen2_0_instruction_master_waitrequest           => nios2_gen2_0_instruction_master_waitrequest,                             --                                           .waitrequest
			nios2_gen2_0_instruction_master_read                  => nios2_gen2_0_instruction_master_read,                                    --                                           .read
			nios2_gen2_0_instruction_master_readdata              => nios2_gen2_0_instruction_master_readdata,                                --                                           .readdata
			hex_digits_pio_s1_address                             => mm_interconnect_0_hex_digits_pio_s1_address,                             --                          hex_digits_pio_s1.address
			hex_digits_pio_s1_write                               => mm_interconnect_0_hex_digits_pio_s1_write,                               --                                           .write
			hex_digits_pio_s1_readdata                            => mm_interconnect_0_hex_digits_pio_s1_readdata,                            --                                           .readdata
			hex_digits_pio_s1_writedata                           => mm_interconnect_0_hex_digits_pio_s1_writedata,                           --                                           .writedata
			hex_digits_pio_s1_chipselect                          => mm_interconnect_0_hex_digits_pio_s1_chipselect,                          --                                           .chipselect
			jtag_uart_0_avalon_jtag_slave_address                 => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address,                 --              jtag_uart_0_avalon_jtag_slave.address
			jtag_uart_0_avalon_jtag_slave_write                   => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write,                   --                                           .write
			jtag_uart_0_avalon_jtag_slave_read                    => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read,                    --                                           .read
			jtag_uart_0_avalon_jtag_slave_readdata                => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata,                --                                           .readdata
			jtag_uart_0_avalon_jtag_slave_writedata               => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata,               --                                           .writedata
			jtag_uart_0_avalon_jtag_slave_waitrequest             => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest,             --                                           .waitrequest
			jtag_uart_0_avalon_jtag_slave_chipselect              => mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect,              --                                           .chipselect
			key_s1_address                                        => mm_interconnect_0_key_s1_address,                                        --                                     key_s1.address
			key_s1_readdata                                       => mm_interconnect_0_key_s1_readdata,                                       --                                           .readdata
			keycode_s1_address                                    => mm_interconnect_0_keycode_s1_address,                                    --                                 keycode_s1.address
			keycode_s1_write                                      => mm_interconnect_0_keycode_s1_write,                                      --                                           .write
			keycode_s1_readdata                                   => mm_interconnect_0_keycode_s1_readdata,                                   --                                           .readdata
			keycode_s1_writedata                                  => mm_interconnect_0_keycode_s1_writedata,                                  --                                           .writedata
			keycode_s1_chipselect                                 => mm_interconnect_0_keycode_s1_chipselect,                                 --                                           .chipselect
			leds_pio_s1_address                                   => mm_interconnect_0_leds_pio_s1_address,                                   --                                leds_pio_s1.address
			leds_pio_s1_write                                     => mm_interconnect_0_leds_pio_s1_write,                                     --                                           .write
			leds_pio_s1_readdata                                  => mm_interconnect_0_leds_pio_s1_readdata,                                  --                                           .readdata
			leds_pio_s1_writedata                                 => mm_interconnect_0_leds_pio_s1_writedata,                                 --                                           .writedata
			leds_pio_s1_chipselect                                => mm_interconnect_0_leds_pio_s1_chipselect,                                --                                           .chipselect
			nios2_gen2_0_debug_mem_slave_address                  => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address,                  --               nios2_gen2_0_debug_mem_slave.address
			nios2_gen2_0_debug_mem_slave_write                    => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write,                    --                                           .write
			nios2_gen2_0_debug_mem_slave_read                     => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read,                     --                                           .read
			nios2_gen2_0_debug_mem_slave_readdata                 => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata,                 --                                           .readdata
			nios2_gen2_0_debug_mem_slave_writedata                => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata,                --                                           .writedata
			nios2_gen2_0_debug_mem_slave_byteenable               => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable,               --                                           .byteenable
			nios2_gen2_0_debug_mem_slave_waitrequest              => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest,              --                                           .waitrequest
			nios2_gen2_0_debug_mem_slave_debugaccess              => mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess,              --                                           .debugaccess
			sdram_s1_address                                      => mm_interconnect_0_sdram_s1_address,                                      --                                   sdram_s1.address
			sdram_s1_write                                        => mm_interconnect_0_sdram_s1_write,                                        --                                           .write
			sdram_s1_read                                         => mm_interconnect_0_sdram_s1_read,                                         --                                           .read
			sdram_s1_readdata                                     => mm_interconnect_0_sdram_s1_readdata,                                     --                                           .readdata
			sdram_s1_writedata                                    => mm_interconnect_0_sdram_s1_writedata,                                    --                                           .writedata
			sdram_s1_byteenable                                   => mm_interconnect_0_sdram_s1_byteenable,                                   --                                           .byteenable
			sdram_s1_readdatavalid                                => mm_interconnect_0_sdram_s1_readdatavalid,                                --                                           .readdatavalid
			sdram_s1_waitrequest                                  => mm_interconnect_0_sdram_s1_waitrequest,                                  --                                           .waitrequest
			sdram_s1_chipselect                                   => mm_interconnect_0_sdram_s1_chipselect,                                   --                                           .chipselect
			sdram_pll_pll_slave_address                           => mm_interconnect_0_sdram_pll_pll_slave_address,                           --                        sdram_pll_pll_slave.address
			sdram_pll_pll_slave_write                             => mm_interconnect_0_sdram_pll_pll_slave_write,                             --                                           .write
			sdram_pll_pll_slave_read                              => mm_interconnect_0_sdram_pll_pll_slave_read,                              --                                           .read
			sdram_pll_pll_slave_readdata                          => mm_interconnect_0_sdram_pll_pll_slave_readdata,                          --                                           .readdata
			sdram_pll_pll_slave_writedata                         => mm_interconnect_0_sdram_pll_pll_slave_writedata,                         --                                           .writedata
			spi_0_spi_control_port_address                        => mm_interconnect_0_spi_0_spi_control_port_address,                        --                     spi_0_spi_control_port.address
			spi_0_spi_control_port_write                          => mm_interconnect_0_spi_0_spi_control_port_write,                          --                                           .write
			spi_0_spi_control_port_read                           => mm_interconnect_0_spi_0_spi_control_port_read,                           --                                           .read
			spi_0_spi_control_port_readdata                       => mm_interconnect_0_spi_0_spi_control_port_readdata,                       --                                           .readdata
			spi_0_spi_control_port_writedata                      => mm_interconnect_0_spi_0_spi_control_port_writedata,                      --                                           .writedata
			spi_0_spi_control_port_chipselect                     => mm_interconnect_0_spi_0_spi_control_port_chipselect,                     --                                           .chipselect
			sysid_qsys_0_control_slave_address                    => mm_interconnect_0_sysid_qsys_0_control_slave_address,                    --                 sysid_qsys_0_control_slave.address
			sysid_qsys_0_control_slave_readdata                   => mm_interconnect_0_sysid_qsys_0_control_slave_readdata,                   --                                           .readdata
			timer_0_s1_address                                    => mm_interconnect_0_timer_0_s1_address,                                    --                                 timer_0_s1.address
			timer_0_s1_write                                      => mm_interconnect_0_timer_0_s1_write,                                      --                                           .write
			timer_0_s1_readdata                                   => mm_interconnect_0_timer_0_s1_readdata,                                   --                                           .readdata
			timer_0_s1_writedata                                  => mm_interconnect_0_timer_0_s1_writedata,                                  --                                           .writedata
			timer_0_s1_chipselect                                 => mm_interconnect_0_timer_0_s1_chipselect,                                 --                                           .chipselect
			usb_gpx_s1_address                                    => mm_interconnect_0_usb_gpx_s1_address,                                    --                                 usb_gpx_s1.address
			usb_gpx_s1_readdata                                   => mm_interconnect_0_usb_gpx_s1_readdata,                                   --                                           .readdata
			usb_irq_s1_address                                    => mm_interconnect_0_usb_irq_s1_address,                                    --                                 usb_irq_s1.address
			usb_irq_s1_readdata                                   => mm_interconnect_0_usb_irq_s1_readdata,                                   --                                           .readdata
			usb_rst_s1_address                                    => mm_interconnect_0_usb_rst_s1_address,                                    --                                 usb_rst_s1.address
			usb_rst_s1_write                                      => mm_interconnect_0_usb_rst_s1_write,                                      --                                           .write
			usb_rst_s1_readdata                                   => mm_interconnect_0_usb_rst_s1_readdata,                                   --                                           .readdata
			usb_rst_s1_writedata                                  => mm_interconnect_0_usb_rst_s1_writedata,                                  --                                           .writedata
			usb_rst_s1_chipselect                                 => mm_interconnect_0_usb_rst_s1_chipselect,                                 --                                           .chipselect
			VGA_text_mode_controller_0_avalon_mm_slave_address    => mm_interconnect_0_vga_text_mode_controller_0_avalon_mm_slave_address,    -- VGA_text_mode_controller_0_avalon_mm_slave.address
			VGA_text_mode_controller_0_avalon_mm_slave_write      => mm_interconnect_0_vga_text_mode_controller_0_avalon_mm_slave_write,      --                                           .write
			VGA_text_mode_controller_0_avalon_mm_slave_read       => mm_interconnect_0_vga_text_mode_controller_0_avalon_mm_slave_read,       --                                           .read
			VGA_text_mode_controller_0_avalon_mm_slave_readdata   => mm_interconnect_0_vga_text_mode_controller_0_avalon_mm_slave_readdata,   --                                           .readdata
			VGA_text_mode_controller_0_avalon_mm_slave_writedata  => mm_interconnect_0_vga_text_mode_controller_0_avalon_mm_slave_writedata,  --                                           .writedata
			VGA_text_mode_controller_0_avalon_mm_slave_byteenable => mm_interconnect_0_vga_text_mode_controller_0_avalon_mm_slave_byteenable, --                                           .byteenable
			VGA_text_mode_controller_0_avalon_mm_slave_chipselect => mm_interconnect_0_vga_text_mode_controller_0_avalon_mm_slave_chipselect  --                                           .chipselect
		);

	irq_mapper : component finalproject_irq_mapper
		port map (
			clk           => clk_clk,                        --       clk.clk
			reset         => rst_controller_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,       -- receiver0.irq
			receiver1_irq => irq_mapper_receiver1_irq,       -- receiver1.irq
			receiver2_irq => irq_mapper_receiver2_irq,       -- receiver2.irq
			sender_irq    => nios2_gen2_0_irq_irq            --    sender.irq
		);

	rst_controller : component finalproject_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,                -- reset_in0.reset
			reset_in1      => nios2_gen2_0_debug_reset_request_reset, -- reset_in1.reset
			clk            => clk_clk,                                --       clk.clk
			reset_out      => rst_controller_reset_out_reset,         -- reset_out.reset
			reset_req      => rst_controller_reset_out_reset_req,     --          .reset_req
			reset_req_in0  => '0',                                    -- (terminated)
			reset_req_in1  => '0',                                    -- (terminated)
			reset_in2      => '0',                                    -- (terminated)
			reset_req_in2  => '0',                                    -- (terminated)
			reset_in3      => '0',                                    -- (terminated)
			reset_req_in3  => '0',                                    -- (terminated)
			reset_in4      => '0',                                    -- (terminated)
			reset_req_in4  => '0',                                    -- (terminated)
			reset_in5      => '0',                                    -- (terminated)
			reset_req_in5  => '0',                                    -- (terminated)
			reset_in6      => '0',                                    -- (terminated)
			reset_req_in6  => '0',                                    -- (terminated)
			reset_in7      => '0',                                    -- (terminated)
			reset_req_in7  => '0',                                    -- (terminated)
			reset_in8      => '0',                                    -- (terminated)
			reset_req_in8  => '0',                                    -- (terminated)
			reset_in9      => '0',                                    -- (terminated)
			reset_req_in9  => '0',                                    -- (terminated)
			reset_in10     => '0',                                    -- (terminated)
			reset_req_in10 => '0',                                    -- (terminated)
			reset_in11     => '0',                                    -- (terminated)
			reset_req_in11 => '0',                                    -- (terminated)
			reset_in12     => '0',                                    -- (terminated)
			reset_req_in12 => '0',                                    -- (terminated)
			reset_in13     => '0',                                    -- (terminated)
			reset_req_in13 => '0',                                    -- (terminated)
			reset_in14     => '0',                                    -- (terminated)
			reset_req_in14 => '0',                                    -- (terminated)
			reset_in15     => '0',                                    -- (terminated)
			reset_req_in15 => '0'                                     -- (terminated)
		);

	rst_controller_001 : component finalproject_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,                -- reset_in0.reset
			reset_in1      => nios2_gen2_0_debug_reset_request_reset, -- reset_in1.reset
			clk            => sdram_pll_c0_clk,                       --       clk.clk
			reset_out      => rst_controller_001_reset_out_reset,     -- reset_out.reset
			reset_req      => open,                                   -- (terminated)
			reset_req_in0  => '0',                                    -- (terminated)
			reset_req_in1  => '0',                                    -- (terminated)
			reset_in2      => '0',                                    -- (terminated)
			reset_req_in2  => '0',                                    -- (terminated)
			reset_in3      => '0',                                    -- (terminated)
			reset_req_in3  => '0',                                    -- (terminated)
			reset_in4      => '0',                                    -- (terminated)
			reset_req_in4  => '0',                                    -- (terminated)
			reset_in5      => '0',                                    -- (terminated)
			reset_req_in5  => '0',                                    -- (terminated)
			reset_in6      => '0',                                    -- (terminated)
			reset_req_in6  => '0',                                    -- (terminated)
			reset_in7      => '0',                                    -- (terminated)
			reset_req_in7  => '0',                                    -- (terminated)
			reset_in8      => '0',                                    -- (terminated)
			reset_req_in8  => '0',                                    -- (terminated)
			reset_in9      => '0',                                    -- (terminated)
			reset_req_in9  => '0',                                    -- (terminated)
			reset_in10     => '0',                                    -- (terminated)
			reset_req_in10 => '0',                                    -- (terminated)
			reset_in11     => '0',                                    -- (terminated)
			reset_req_in11 => '0',                                    -- (terminated)
			reset_in12     => '0',                                    -- (terminated)
			reset_req_in12 => '0',                                    -- (terminated)
			reset_in13     => '0',                                    -- (terminated)
			reset_req_in13 => '0',                                    -- (terminated)
			reset_in14     => '0',                                    -- (terminated)
			reset_req_in14 => '0',                                    -- (terminated)
			reset_in15     => '0',                                    -- (terminated)
			reset_req_in15 => '0'                                     -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;

	mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;

	mm_interconnect_0_sdram_s1_read_ports_inv <= not mm_interconnect_0_sdram_s1_read;

	mm_interconnect_0_sdram_s1_byteenable_ports_inv <= not mm_interconnect_0_sdram_s1_byteenable;

	mm_interconnect_0_sdram_s1_write_ports_inv <= not mm_interconnect_0_sdram_s1_write;

	mm_interconnect_0_keycode_s1_write_ports_inv <= not mm_interconnect_0_keycode_s1_write;

	mm_interconnect_0_usb_rst_s1_write_ports_inv <= not mm_interconnect_0_usb_rst_s1_write;

	mm_interconnect_0_hex_digits_pio_s1_write_ports_inv <= not mm_interconnect_0_hex_digits_pio_s1_write;

	mm_interconnect_0_leds_pio_s1_write_ports_inv <= not mm_interconnect_0_leds_pio_s1_write;

	mm_interconnect_0_timer_0_s1_write_ports_inv <= not mm_interconnect_0_timer_0_s1_write;

	mm_interconnect_0_spi_0_spi_control_port_read_ports_inv <= not mm_interconnect_0_spi_0_spi_control_port_read;

	mm_interconnect_0_spi_0_spi_control_port_write_ports_inv <= not mm_interconnect_0_spi_0_spi_control_port_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

	rst_controller_001_reset_out_reset_ports_inv <= not rst_controller_001_reset_out_reset;

end architecture rtl; -- of finalproject
